000|T121|5-FU
000|T121|leucovorin
000|T121|oxaliplatin
000|T121|FOLFOX 6