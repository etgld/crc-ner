0|today
0|ate
0|ton
0|TON
0|yesterday
0|thursday
0|friday
0|january