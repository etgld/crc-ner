000|T121|cytoxan
000|T121|taxotere
000|T121|tamoxifen
000|T121|chemotherapy
000|T121|TC
000|T121|chemo