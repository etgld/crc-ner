000|T121|TC
000|T121|cisplatin
000|T121|gemcitabine
000|T121|Doxcil
000|T121|Carboplatin
000|T121|Taxol