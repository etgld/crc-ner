T051|today
T051|ate
T051|ton
T051|TON
T051|yesterday
T051|thursday
T051|friday
T051|january
T051|5