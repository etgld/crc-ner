000|T121|chemotherapy
000|T121|chemotherapies
000|T121|chemo
000|T121|chemotherapeutic
000|T121|liposomal doxorubicin
000|T121|carboplatin
000|T121|paclitaxel
000|T121|gemcitabine
000|T121|cisplatin
000|T121|platinum
000|T121|doxil
000|T121|taxol
000|T121|ataxol
000|T121|carbo
000|T121|gemzar
000|T121|topotecan
000|T121|carbotaxol