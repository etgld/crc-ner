000|T121|-20-2011
000|T121|.
000|T121|. if neoadj
000|T121|. she
000|T121|01-29-2002
000|T121|01230 reco
000|T121|09-24-2010
000|T121|10118 re
000|T121|10930 re
000|T121|1112 recor
000|T121|20314 reco
000|T121|20403 reco
000|T121|20801 reco
000|T121|20815 reco
000|T121|21128 reco
000|T121|30816 re
000|T121|31001 reco
000|T121|31008 reco
000|T121|4fu
000|T121|5-f
000|T121|5-fluorouracil
000|T121|5-fu
000|T121|5f-u
000|T121|5fu
000|T121|6-mp
000|T121|a testin
000|T121|a.c
000|T121|a/c
000|T121|about was t
000|T121|abraxan
000|T121|abraxane
000|T121|abvd
000|T121|ac
000|T121|ac-t
000|T121|act
000|T121|adalimumab
000|T121|adriamy
000|T121|adriamycin
000|T121|adrucil
000|T121|afiblercept
000|T121|aflibercept
000|T121|alfa-2b interferon
000|T121|alflibercept
000|T121|alibercept
000|T121|alpha 2b interferon
000|T121|alpha interferon
000|T121|alpha-2b interferon
000|T121|an oncotype
000|T121|anastrazole
000|T121|anastrozole
000|T121|and her fam
000|T121|anthracycline
000|T121|arimedex
000|T121|arimidex
000|T121|aromasin
000|T121|aromatase
000|T121|aromatase inhibitor
000|T121|as breast c
000|T121|as diff
000|T121|ase a
000|T121|ataxol
000|T121|ativan
000|T121|avastin
000|T121|avstin
000|T121|aware
000|T121|azathioprine
000|T121|bev
000|T121|bevacizumab
000|T121|bolus 5-fu
000|T121|bout a 20% c
000|T121|caboplatin
000|T121|cabotaxol
000|T121|capecitabine
000|T121|capeox
000|T121|capptosar
000|T121|carbo
000|T121|carbo-taxol
000|T121|carboplat
000|T121|carboplatin
000|T121|carboplatinum
000|T121|carbotaxol
000|T121|cetuximab
000|T121|chem
000|T121|chemo
000|T121|chemo radiation
000|T121|chemo therapy
000|T121|chemo-radiation
000|T121|chemo-rt
000|T121|chemoembolization
000|T121|chemoirradiation
000|T121|chemorad
000|T121|chemoradiation
000|T121|chemoradiotherapy
000|T121|chemort
000|T121|chemotherap
000|T121|chemotherapeutic
000|T121|chemotherapies
000|T121|chemotherapy
000|T121|chemotherapy's
000|T121|chemotheray
000|T121|chmeo
000|T121|cisplatin
000|T121|cistoplatin
000|T121|cpt-11
000|T121|cyclophosphamide
000|T121|cytotaxin
000|T121|cytoxan
000|T121|cytoxan pr
000|T121|d cytoxan.
000|T121|d have very
000|T121|dalotuzumab
000|T121|denies
000|T121|denosumab
000|T121|docetaxel
000|T121|docetaxil
000|T121|docetaxol
000|T121|doxil
000|T121|doxorubicin
000|T121|e gaining iv
000|T121|ection with
000|T121|ed in deta
000|T121|ed plan. s
000|T121|edical histo
000|T121|eloxatin
000|T121|ent due to t
000|T121|erbitux
000|T121|ery well
000|T121|etoposide
000|T121|examestane
000|T121|exemestane
000|T121|femara
000|T121|fluorburacil
000|T121|fluoropyrimidine
000|T121|fluorouracil
000|T121|folferi
000|T121|folfiri
000|T121|folfirinox
000|T121|folfox
000|T121|folfox 6
000|T121|folfox 7
000|T121|folfox therapy
000|T121|folfox-6
000|T121|folfox-iri
000|T121|folfox6
000|T121|folfox7
000|T121|folfoxiri
000|T121|for 2 w
000|T121|for 5
000|T121|for breast
000|T121|fulvestrant
000|T121|gemcitabine
000|T121|gemzar
000|T121|he is being
000|T121|he is i
000|T121|herapy and
000|T121|herceptin
000|T121|hipec
000|T121|humira
000|T121|i-131
000|T121|id recommend
000|T121|ihcp
000|T121|il 2
000|T121|il-2
000|T121|il2
000|T121|in det
000|T121|in the prim
000|T121|infliximab
000|T121|inteferon
000|T121|interferon
000|T121|interferon, alpha 2b
000|T121|interleukin
000|T121|interleukin 2
000|T121|interleukin-2
000|T121|intraperitoneal hyperthemic chemoperfusion
000|T121|ipilimumab
000|T121|irection of
000|T121|irinotecan
000|T121|is er posit
000|T121|is not compl
000|T121|ively as her
000|T121|l allow us t
000|T121|l risks, b
000|T121|leucovorin
000|T121|liposomal doxorubicin
000|T121|lonsurf
000|T121|lupron
000|T121|maid
000|T121|melphalan
000|T121|ment sche
000|T121|mercaptopurine
000|T121|methotrexate
000|T121|mfolfox 6
000|T121|mfolfox-6
000|T121|mfolfox6
000|T121|mitomycin
000|T121|mitomycin c
000|T121|mitomycin-c
000|T121|mopp
000|T121|n and ar
000|T121|nce of progr
000|T121|neulasta
000|T121|nse of the t
000|T121|ntact
000|T121|oceeding wit
000|T121|of concerni
000|T121|of the brai
000|T121|on186, ph
000|T121|or to breast
000|T121|otherapy. i
000|T121|oughout her
000|T121|ould like to
000|T121|oxali
000|T121|oxaliplatin
000|T121|oxalplatin
000|T121|oxaplatin
000|T121|paciltaxel
000|T121|paclitaxel
000|T121|paclitaxela
000|T121|panitumumab
000|T121|paraplatin
000|T121|patient was
000|T121|paxil
000|T121|perjeta
000|T121|platinum
000|T121|post
000|T121|prechemotherapy
000|T121|radiochemotherapy
000|T121|rapy. pathol
000|T121|regorafenib
000|T121|remicade
000|T121|ridafololimus
000|T121|ridosol
000|T121|ritux
000|T121|rituximab
000|T121|rson132, d
000|T121|s therapy
000|T121|seen person
000|T121|she is curre
000|T121|she stat
000|T121|sorafenib
000|T121|stions,
000|T121|t/c
000|T121|tamoxifen
000|T121|tasisulam
000|T121|tax
000|T121|taxane
000|T121|taxo
000|T121|taxol
000|T121|taxotere
000|T121|taxtotere
000|T121|tc
000|T121|tch
000|T121|temozolomide
000|T121|tient st
000|T121|today. we w
000|T121|topotecan
000|T121|toxicity
000|T121|ts, and
000|T121|vaccinia
000|T121|vaccinia virus
000|T121|vectibix
000|T121|vomiting, es
000|T121|was stop
000|T121|were ans
000|T121|x 1 year
000|T121|x 5 year
000|T121|xeliri
000|T121|xeloda
000|T121|xelox
000|T121|xgeva
000|T121|y problems
000|T121|zometa