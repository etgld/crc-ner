00000|T121|Capecitabine monotherapy
00000|T121|Capecitabine (Xeloda)
00000|T121|Oxaliplatin (Eloxatin)
00000|T121|Fluorouracil (5-FU)
00000|T121|Folinic acid (Leucovorin)
00000|T121|Levoleucovorin (Fusilev)
00000|T121|Tegafur and uracil (UFT)
00000|T121|Irinotecan (Camptosar)
00000|T121|Floxuridine (FUDR)
00000|T121|Mitomycin (Mutamycin)
00000|T121|Trifluridine and tipiracil (Lonsurf)
00000|T121|Trifluridine and tipiracil monotherapy
00000|T121|Irinotecan monotherapy
00000|T121|FULV & Bevacizumab
00000|T121|FOLFOX4 & Bevacizumab
00000|T121|FOLFOX4 (L-Leucovorin)
00000|T121|FOLFOX4
00000|T121|Fluorouracil monotherapy
00000|T121|FOLFIRI
00000|T121|CapeOx (XELOX)
00000|T121|IROX
00000|T121|IRIS
00000|T121|mFOLFOX6-B
00000|T121|mFOLFOX6
00000|T121|FOLFIRI & Ziv-aflibercept
00000|T121|FOLFIRI & Ramucirumab
00000|T121|FOLFIRI & Bevacizumab
00000|T121|FOLFIRI (L-Leucovorin)
00000|T121|CAPIRI-Bev
00000|T121|CAPIRI
00000|T121|CapeIRI
00000|T121|mXELIRI & Bevacizumab
00000|T121|CAPIRI
00000|T121|XELIRI
00000|T121|mXELIRI
00000|T121|CapeOx & Erlotinib
00000|T121|XELOX
00000|T121|S-1 monotherapy
00000|T121|Fluorouracil & Bevacizumab
00000|T121|Tegafur, gimeracil, oteracil (S-1)
00000|T121|SOX & Bevacizumab
00000|T121|OXAFAFU
00000|T121|Nordic FLOX
00000|T121|IFL
00000|T121|mIFL
00000|T121|FUOX
00000|T121|FULV (L-Leucovorin)
00000|T121|FULV
00000|T121|FUIRI
00000|T121|mFOLFOX6-B (L-Leucovorin)
00000|T121|mFOLFOX6-B
00000|T121|FOLFOX-B
00000|T121|mFOLFOX7
00000|T121|mFOLFOX7 (L-Leucovorin)
00000|T121|FOLFOX 7/sLV5FU2 (L-Leucovorin)
00000|T121|FOLFOX 7/sLV5FU2
00000|T121|mFOLFOX6 (L-Leucovorin)
00000|T121|FOLFOX2
00000|T121|FOLFIRINOX & Bevacizumab (L-Leucovorin)
00000|T121|FOLFIRINOX & Bevacizumab
00000|T121|FOLFOXIRI & Bevacizumab
00000|T121|FOLFIRINOX
00000|T121|FOLFOXIRI
00000|T121|FOLFIRI & Bevacizumab (L-Leucovorin)
00000|T121|CAPIRI-Bev
00000|T121|XELIRI-Bev
00000|T121|CapeOx & Bevacizumab
00000|T121|CAPOX-B
00000|T121|XELOX & Bevacizumab
00000|T121|COX
00000|T121|Capecitabine & Bevacizumab
00000|T121|Tegafur, Uracil, Folinic acid
00000|T121|Tegafur and uracil (UFT)
00000|T121|UFT + LV
