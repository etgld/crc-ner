35802855|T121|AMG 330
35802856|T121|AZD5363
35802856|T121|Capivasertib
35802857|T121|Abciximab
35802858|T121|LY2835219
35802858|T121|Abemaciclib
35802859|T121|PCI-24781
35802859|T121|Abexinostat
35802860|T121|CB7630
35802860|T121|abiraterone acetate
35802860|T121|Abiraterone
35802861|T121|ACP-196
35802861|T121|Acalabrutinib
35802862|T121|paracetamol
35802862|T121|paracetamole
35802862|T121|APAP
35802862|T121|Acetaminophen
35802863|T121|MA144-A1
35802863|T121|aclacinomycin
35802863|T121|aclacinomycin A hydrochloride
35802863|T121|aclacinomycin-A
35802863|T121|aclarubicin hydrochloride
35802863|T121|aclacinomycin A
35802863|T121|Aclarubicin
35802864|T121|Actinium Ac 225 lintuzumab
35802865|T121|ACV
35802865|T121|acycloguanosine
35802865|T121|aciclovir
35802865|T121|Acyclovir
35802866|T121|ado-trastuzumab emtansine
35802866|T121|Ado-trastuzumab emtansine
35802866|T121|PRO132365
35802866|T121|TDM1
35802866|T121|T-DM1
35802866|T121|Trastuzumab emtansine
35802867|T121|BIBW-2992
35802867|T121|afatinib dimaleate
35802867|T121|BIBW 2992
35802867|T121|Afatinib
35802868|T121|GSK2110183
35802868|T121|Afuresertib
35802869|T121|IL-2
35802869|T121|Interleukin-2
35802869|T121|Aldesleukin
35802870|T121|AF802
35802870|T121|AF-802
35802870|T121|RG7853
35802870|T121|RO5424802
35802870|T121|UNII-LIJ4CT1Z3Y
35802870|T121|CH5424802
35802870|T121|Alectinib
35802871|T121|LDP03
35802871|T121|Alemtuzumab
35802872|T121|acido alendronico
35802872|T121|alendronic acid
35802872|T121|acide alendronique
35802872|T121|Alendronate
35802873|T121|MLN8237
35802873|T121|Alisertib
35802874|T121|all-trans retinoic acid
35802874|T121|ATRA
35802874|T121|tretinoin
35802874|T121|All-trans retinoic acid
35802875|T121|Allopurinol
35802876|T121|Alprazolam
35802877|T121|hexamethylmelamine
35802877|T121|HMM
35802877|T121|Altretamine
35802878|T121|L-868275
35802878|T121|flavopiridol
35802878|T121|HMR 1275
35802878|T121|Alvocidib
35802879|T121|MORAb-009
35802879|T121|Amatuximab
35802880|T121|Amifostine
35802881|T121|6-aminohexanoic acid
35802881|T121|ε-aminocaproic acid
35802881|T121|ε-Ahx
35802881|T121|epsilon aminocaproic acid
35802881|T121|Aminocaproic acid
35802882|T121|Aminoglutethimide
35802883|T121|Aminopterin
35802884|T121|SM-5887
35802884|T121|AMR
35802884|T121|amrubicin HCI
35802884|T121|Amrubicin
35802885|T121|SN-11841
35802885|T121|acridinyl anisidide
35802885|T121|AMSA
35802885|T121|Cain's acridine
35802885|T121|m-AMSA
35802885|T121|CI-880
35802885|T121|Amsacrine
35802886|T121|Anagrelide
35802887|T121|Anastrozole
35802888|T121|Anti-inhibitor coagulant complex
35802889|T121|Antithrombin III
35802890|T121|Antithymocyte globulin horse ATG
35802891|T121|anti-thymocyte globulin (rabbit)
35802891|T121|lymphocyte immune globulin (rabbit)
35802891|T121|antithymocyte globulin (rabbit)
35802891|T121|Antithymocyte globulin rabbit ATG
35802892|T121|ARN-509
35802892|T121|Apalutamide
35802893|T121|YN968D1
35802893|T121|rivoceranib
35802893|T121|Apatinib
35802894|T121|Apixaban
35802895|T121|MK-0869
35802895|T121|Aprepitant
35802896|T121|Argatroban
35802897|T121|Arsenic trioxide
35802898|T121|colaspase
35802898|T121|L Asparaginase
35802898|T121|L-ASP
35802898|T121|crisantaspase
35802898|T121|Asparaginase
35802899|T121|crisantaspasum
35802899|T121|crisantaspase
35802899|T121|krisantaspaasi
35802899|T121|krisantaspas
35802899|T121|Erwinia L-asparginase
35802899|T121|Asparaginase Erwinia chrysanthemi
35802900|T121|A.A.S.
35802900|T121|A.S.A.
35802900|T121|AAC
35802900|T121|AAS
35802900|T121|Acetylsalicylate Calcium
35802900|T121|Acetylsalicylate Copper
35802900|T121|Acetylsalicylate Lysine
35802900|T121|Acetylsalicylate Sodium
35802900|T121|Acetylsalicylic Acid Aluminium
35802900|T121|Acetylsalicylic Acid Effervescent
35802900|T121|Acetylsalicylic Acid Enteric Coated
35802900|T121|Acid Acetylsalicylic
35802900|T121|A-A-S 500
35802900|T121|Acidum Acethylsalicylicum
35802900|T121|Acidum Acetylsalicum
35802900|T121|Acidum Acetylsalicylic
35802900|T121|Acidum Acetylsalicylicum
35802900|T121|Acidum Ascorbinicum
35802900|T121|ASA
35802900|T121|ASS
35802900|T121|ECASA
35802900|T121|Methyl Diethylacetylsalicylate
35802900|T121|Aspirin
35802900|T121|Acido Acetilsalicilico
35802901|T121|Aspirin and dipyridamole
35802902|T121|MPDL3280A
35802902|T121|RG7446
35802902|T121|RO5541267
35802902|T121|Atezolizumab
35802903|T121|Atovaquone
35802904|T121|Atropine
35802905|T121|YM477
35802905|T121|AKR 501
35802905|T121|E5501
35802905|T121|Avatrombopag
35802906|T121|MSB0010718C
35802906|T121|Avelumab
35802907|T121|Axicel
35802907|T121|Axi-cel
35802907|T121|KTE-C19
35802907|T121|Axicabtagene ciloleucel
35802908|T121|AG013736
35802908|T121|AG-013736
35802908|T121|Axitinib
35802909|T121|5-azacitidine
35802909|T121|5-azacytidine
35802909|T121|Azacitidine
35802910|T121|BHQ880
35802911|T121|GCR-3888
35802911|T121|CAT-3888
35802911|T121|BL22 immunotoxin
35802912|T121|Bacille Calmette–Guerin
35802912|T121|Bacillus Calmette-Guerin
35802913|T121|AZD1152
35802913|T121|Barasertib
35802914|T121|PGN401
35802914|T121|Bavituximab
35802915|T121|Belagenpumatucel-L
35802916|T121|PXD101
35802916|T121|Belinostat
35802917|T121|CKD-602
35802917|T121|belotecan hydrochloride
35802917|T121|Belotecan
35802918|T121|CEP-18083
35802918|T121|SDX-105
35802918|T121|SyB L-0501
35802918|T121|bendamustine hydrochloride
35802918|T121|cytostasan hydrochloride
35802918|T121|bendamustin hydrochloride
35802918|T121|Bendamustine
35802919|T121|PRT-054021
35802919|T121|Betrixaban
35802920|T121|ABP 215
35802920|T121|Bevacizumab-awwb
35802921|T121|rhuMab-VEGF
35802921|T121|Bevacizumab
35802922|T121|LGD1069
35802922|T121|Bexarotene
35802923|T121|Bicalutamide
35802924|T121|ARRY-162
35802924|T121|ARRY-438162
35802924|T121|MEK162
35802924|T121|Binimetinib
35802925|T121|Bivalirudin
35802926|T121|Bleomycin
35802927|T121|AMG 103
35802927|T121|MEDI538
35802927|T121|MT103
35802927|T121|Blinatumomab
35802928|T121|MLN341
35802928|T121|PS-341
35802928|T121|LDP 341
35802928|T121|Bortezomib
35802929|T121|SKI-606
35802929|T121|Bosutinib
35802930|T121|cAC10-vcMMAE
35802930|T121|SGN-35
35802930|T121|Brentuximab vedotin
35802931|T121|AP26113
35802931|T121|Brigatinib
35802932|T121|BKM120
35802932|T121|Buparlisib
35802933|T121|Busulfan
35802934|T121|XRP6258
35802934|T121|TXD258
35802934|T121|RPR116258A
35802934|T121|Cabazitaxel
35802935|T121|XL-184
35802935|T121|XL184
35802935|T121|Cabozantinib
35802936|T121|calaspargase pegol-mknl
35802936|T121|Calaspargase
35802937|T121|artificial saliva
35802937|T121|supersaturated calcium phosphate rinse
35802937|T121|Calcium phosphate rinse
35802938|T121|Cangrelor
35802939|T121|Ro 09-1978/000
35802939|T121|capecitabine RDT
35802939|T121|kapesitabin
35802939|T121|Capecitabine
35802940|T121|ALX-0081
35802940|T121|caplacizumab-yhdp
35802940|T121|Caplacizumab
35802941|T121|JM8
35802941|T121|Carboplatin
35802942|T121|CFZ
35802942|T121|PR-171
35802942|T121|Carfilzomib
35802943|T121|BCNU
35802943|T121|bischloroethylnitrosourea
35802943|T121|carmustin
35802943|T121|Carmustine
35802944|T121|NPC-08
35802944|T121|NSC-409962
35802944|T121|WR-139021
35802944|T121|polifeprosan 20 with carmustine implant
35802944|T121|Carmustine wafer polifeprosan 20
35802945|T121|Caspofungin
35802946|T121|Catumaxomab
35802947|T121|AZD2171
35802947|T121|Cediranib
35802948|T121|REGN2810
35802948|T121|cemiplimab-rwlc
35802948|T121|Cemiplimab
35802949|T121|LDK378
35802949|T121|Ceritinib
35802950|T121|Cetirizine
35802951|T121|C225
35802951|T121|Cetuximab
35802952|T121|CS055
35802952|T121|HBI-8000
35802952|T121|tucidinostat
35802952|T121|Chidamide
35802953|T121|Chlorambucil
35802954|T121|chlorphenamine
35802954|T121|Chlorpheniramine
35802955|T121|Cilostazol
35802956|T121|Cimetidine
35802957|T121|Ciprofloxacin
35802958|T121|CDDP
35802958|T121|cis-diamminedichloroplatinum III
35802958|T121|cis-platinum
35802958|T121|NSC 119875
35802958|T121|DACP
35802958|T121|DDP
35802958|T121|cisplatinum
35802958|T121|Cisplatin
35802959|T121|IMC-A12
35802959|T121|Cixutumumab
35802960|T121|2-chlorodeoxyadenosine
35802960|T121|2-CdA
35802960|T121|Cladribine
35802961|T121|Clarithromycin
35802962|T121|Clemastine
35802963|T121|clodronate disodium
35802963|T121|clodronic acid disodium tetrahydrate
35802963|T121|Clodronate
35802964|T121|klofarabin
35802964|T121|Clofarabine
35802965|T121|Clopidogrel
35802966|T121|XL518
35802966|T121|GDC-0973
35802966|T121|Cobimetinib
35802967|T121|SAR3419
35802967|T121|CoR
35802967|T121|Coltuximab ravtansine
35802968|T121|BAY 80-6946
35802968|T121|Copanlisib
35802969|T121|Cortisone
35802970|T121|CP-868-596
35802970|T121|Crenolanib
35802971|T121|crizanlizumab-tmca
35802971|T121|SEG101
35802971|T121|Crizanlizumab
35802972|T121|PF02341066
35802972|T121|PF-02341066
35802972|T121|Crizotinib
35802973|T121|OGX-011
35802973|T121|Custirsen
35802974|T121|cobalamin
35802974|T121|vitamin B12
35802974|T121|vitamin B-12
35802974|T121|Cyanocobalamin
35802975|T121|B-518
35802975|T121|WR-138719
35802975|T121|CP monohydrate
35802975|T121|Asta B 518
35802975|T121|cyclophosphamid monohydrate
35802975|T121|cyclophosphamide monohydrate
35802975|T121|CPM
35802975|T121|Cyclophosphamide
35802976|T121|Cyclosporine modified
35802977|T121|Cyclosporine non-modified
35802978|T121|Cyproterone acetate
35802979|T121|Ara-C
35802979|T121|arabinofuranosyl cytidine
35802979|T121|cytosine arabinoside
35802979|T121|arabinosylcytosine
35802979|T121|Cytarabine
35802980|T121|CPX-351
35802980|T121|Cytarabine and daunorubicin liposomal
35802981|T121|Liposomal Ara-C
35802981|T121|Cytarabine liposomal
35802982|T121|Cytomegalovirus Immune Globulin
35802983|T121|Dabigatran
35802984|T121|GSK-2118436A
35802984|T121|dabrafenib mesylate
35802984|T121|GSK2118436
35802984|T121|Dabrafenib
35802985|T121|dacarbazin
35802985|T121|imidazole carboxamide
35802985|T121|DTIC
35802985|T121|Dacarbazine
35802986|T121|PF-00299804
35802986|T121|Dacomitinib
35802987|T121|AC-DE
35802987|T121|actinomycin D
35802987|T121|Dactinomycin
35802988|T121|Dalteparin
35802989|T121|Danaparoid
35802990|T121|Danazol
35802991|T121|Dapsone
35802992|T121|JNJ-54767414
35802992|T121|daratumumab-fihj
35802992|T121|Daratumumab
35802993|T121|Darbepoetin alfa
35802994|T121|ODM-201
35802994|T121|BAY-1841788
35802994|T121|Darolutamide
35802995|T121|BMS-354825
35802995|T121|Dasatinib
35802996|T121|daunomycin
35802996|T121|Daunorubicin
35802997|T121|daunorubicin citrate liposome injection
35802997|T121|Daunorubicin liposomal
35802998|T121|5-aza-2'-deoxycytidine
35802998|T121|Decitabine
35802999|T121|Deferasirox
35803000|T121|Deferiprone
35803001|T121|desferrioxamine B
35803001|T121|desferoxamine B
35803001|T121|DFOA
35803001|T121|DFB
35803001|T121|DFO-B
35803001|T121|Deferoxamine
35803002|T121|polydeoxyribonucleotide sodium salt
35803002|T121|Defibrotide
35803003|T121|FE200486
35803003|T121|degarelix acetate
35803003|T121|ASP3550
35803003|T121|Degarelix
35803004|T121|DAB(389)-interleukin-2
35803004|T121|DAB389 interleukin-2
35803004|T121|DABIL2
35803004|T121|LY335348
35803004|T121|DAB389 interleukin-2 immunotoxin
35803004|T121|Denileukin diftitox
35803005|T121|SGN-CD19A
35803005|T121|Denintuzumab mafodotin
35803006|T121|Denosumab
35803007|T121|Desmopressin
35803008|T121|dexamethasone sodium
35803008|T121|dexamethasone sodium metasulfobenzoate
35803008|T121|dexamethasone sodium phosphate
35803008|T121|dexamethasone acetate
35803008|T121|dexamethasone sodium sulfate
35803008|T121|dexamethasone sodium succinate
35803008|T121|Dexamethasone
35803009|T121|Dexchlorpheniramine
35803010|T121|ADR-529
35803010|T121|ICRF-187
35803010|T121|dexrazoxane hydrochloride
35803010|T121|Dexrazoxane
35803011|T121|stilbestrol
35803011|T121|stilboestrol
35803011|T121|DES
35803011|T121|Diethylstilbestrol
35803012|T121|MK-7965
35803012|T121|SCH 727965
35803012|T121|Dinaciclib
35803013|T121|Ch14.18
35803013|T121|MOAB Ch14.18
35803013|T121|monoclonal antibody Ch14.18
35803013|T121|Dinutuximab
35803014|T121|Diphenhydramine
35803015|T121|Dipyridamole
35803016|T121|RP 56976
35803016|T121|NSC 628503
35803016|T121|Docetaxel
35803017|T121|Docusate
35803018|T121|dolasetron mesylate
35803018|T121|Dolasetron
35803019|T121|Domperidone
35803020|T121|CHIR-258
35803020|T121|TKI-258
35803020|T121|Dovitinib lactate
35803020|T121|Dovitinib
35803021|T121|Doxifluridine
35803022|T121|FI-106
35803022|T121|ADM
35803022|T121|doxorubicin hydrochloride
35803022|T121|hydroxydaunorubicin
35803022|T121|Doxorubicin
35803023|T121|Doxycycline
35803024|T121|Dronabinol
35803025|T121|MEDI4736
35803025|T121|Durvalumab
35803026|T121|Dutasteride
35803027|T121|IPI-145
35803027|T121|Duvelisib
35803028|T121|Eculizumab
35803029|T121|DU-176b
35803029|T121|Edoxaban
35803030|T121|Edrecolomab
35803031|T121|HuLuc63
35803031|T121|PDL063
35803031|T121|PDL-063
35803031|T121|anti-CS1 monoclonal antibody HuLuc63
35803031|T121|BMS-901608
35803031|T121|Elotuzumab
35803032|T121|SB-497115-GR
35803032|T121|Eltrombopag
35803033|T121|ACE910
35803033|T121|emicizumab-kxwh
35803033|T121|Emicizumab
35803034|T121|AG-221
35803034|T121|CC-90007
35803034|T121|enasidenib mesylate
35803034|T121|Enasidenib
35803035|T121|LGX818
35803035|T121|Encorafenib
35803036|T121|Enoxaparin
35803037|T121|X-396
35803037|T121|Ensartinib
35803038|T121|MS-275
35803038|T121|SNDX-275
35803038|T121|Entinostat
35803039|T121|GS-9973
35803039|T121|Entospletinib
35803040|T121|RXDX-101
35803040|T121|Entrectinib
35803041|T121|MDV3100
35803041|T121|Enzalutamide
35803042|T121|Epinephrine autoinjector
35803043|T121|4-epi-doxorubicin
35803043|T121|epidoxorubicin
35803043|T121|Epirubicin
35803044|T121|Epoetin alfa-epbx
35803045|T121|Erythropoetin
35803045|T121|Erythropoietin
35803045|T121|Epoetin alfa
35803046|T121|hLL2
35803046|T121|AMG 412
35803046|T121|Epratuzumab
35803047|T121|Eptifibatide
35803048|T121|JNJ-42756493
35803048|T121|Erdafitinib
35803049|T121|E7389
35803049|T121|ER-086526
35803049|T121|eribulin mesylate
35803049|T121|NSC-707389
35803049|T121|Eribulin
35803050|T121|CP-358
35803050|T121|CP-774
35803050|T121|erlotinib hydrochloride
35803050|T121|OSI-774
35803050|T121|Erlotinib
35803051|T121|estradiol valerate
35803051|T121|estrogens conjugated
35803051|T121|estrogens esterified
35803051|T121|Estradiol
35803052|T121|estramustine phosphate sodium
35803052|T121|Estramustine
35803053|T121|VP-16
35803053|T121|VP-TEC
35803053|T121|VP 16213
35803053|T121|etoposide phosphate
35803053|T121|Etoposide
35803054|T121|RAD001
35803054|T121|RAD-001
35803054|T121|Everolimus
35803055|T121|FCE-24304
35803055|T121|Exemestane
35803056|T121|coagulation factor 9
35803056|T121|FIX
35803056|T121|Christmas Factor
35803056|T121|Factor IX human
35803057|T121|recombinant Christmas Factor
35803057|T121|recombinant FIX
35803057|T121|recombinant coagulation factor 9
35803057|T121|Factor IX recombinant
35803058|T121|Factor IX recombinant Fc fusion protein
35803059|T121|coagulation factor 8
35803059|T121|Factor VIII human
35803060|T121|recombinant coagulation factor 8
35803060|T121|Factor VIII recombinant
35803061|T121|recombinant coagulation factor VIIa
35803061|T121|eptacog alfa (activated)
35803061|T121|recombinant factor 7a
35803061|T121|Factor VIIa recombinant
35803062|T121|FXIII
35803062|T121|coagulation factor 13
35803062|T121|Factor XIII concentrate human
35803063|T121|PRT4445
35803063|T121|andexanet alfa
35803063|T121|Factor Xa recombinant inactivated-zhzo
35803064|T121|Famciclovir
35803065|T121|Famotidine
35803066|T121|Ferric carboxymaltose
35803067|T121|sodium ferric gluconate complex in sucrose injection
35803067|T121|Ferric gluconate
35803068|T121|Ferrous sulfate
35803069|T121|Ferumoxytol
35803070|T121|ARRY-520
35803070|T121|Filanesib
35803071|T121|Filgrastim-sndz
35803072|T121|GCSF
35803072|T121|G-CSF
35803072|T121|granulocyte colony stimulating factor
35803072|T121|filgrastim
35803072|T121|Filgrastim
35803073|T121|Finasteride
35803074|T121|floxuridin
35803074|T121|fluorodeoxyuridine
35803074|T121|fluorouridine deoxyribose
35803074|T121|WR-138720
35803074|T121|Floxuridine
35803075|T121|Fluconazole
35803076|T121|fludarabine phosphate
35803076|T121|FAMP
35803076|T121|Fludarabine
35803077|T121|5 Fluorouracil
35803077|T121|5 FU
35803077|T121|5-FU
35803077|T121|5-fluoracilo
35803077|T121|5-fluorouracilo
35803077|T121|5-fluorouracyl
35803077|T121|FU
35803077|T121|Ro-2-9757
35803077|T121|Fluorouracil
35803078|T121|Fluoxymesterone
35803079|T121|Flutamide
35803080|T121|Folic acid
35803081|T121|calcium folinate
35803081|T121|folinate calcium
35803081|T121|folinato de calcio
35803081|T121|leucovorin calcium
35803081|T121|citrovorum factor
35803081|T121|sodium folinate
35803081|T121|LV
35803081|T121|Folinic acid
35803082|T121|Fondaparinux
35803083|T121|Formestane
35803084|T121|BCX-1777
35803084|T121|immucillin H
35803084|T121|Forodesine
35803085|T121|fosaprepitant dimeglumine
35803085|T121|Fosaprepitant
35803086|T121|R935788
35803086|T121|R788
35803086|T121|Fostamatinib
35803087|T121|Fotemustine
35803088|T121|HMPL-013
35803088|T121|Fruquintinib
35803089|T121|ICI 182780
35803089|T121|ZD9238
35803089|T121|Fulvestrant
35803090|T121|Furosemide
35803091|T121|AR-V7
35803091|T121|TOK-001
35803091|T121|VN/124-1
35803091|T121|Galeterone
35803092|T121|STA-9090
35803092|T121|Ganetespib
35803093|T121|AMG 479
35803093|T121|Ganitumab
35803094|T121|ZD1839
35803094|T121|Gefitinib
35803095|T121|LY-188011
35803095|T121|difluorodeoxycytidine hydrochloride
35803095|T121|gemcitabine hydrochloride
35803095|T121|Gemcitabine
35803096|T121|Gemtuzumab ozogamicin
35803097|T121|ASP2215
35803097|T121|Gilteritinib
35803098|T121|PF-04449913
35803098|T121|Glasdegib
35803099|T121|carboxypeptidase G2
35803099|T121|Glucarpidase
35803100|T121|goserelin acetate
35803100|T121|Goserelin
35803101|T121|granisetron extended-release injection for subcutaneous use
35803101|T121|granisetron hydrochloride
35803101|T121|granisetron hydroxychloride extended release
35803101|T121|granisetron transdermal system
35803101|T121|granisetronum
35803101|T121|Granisetron
35803102|T121|SGI-110
35803102|T121|S110
35803102|T121|Guadecitabine
35803103|T121|Haloperidol
35803104|T121|Hematopoetic progenitor cells cord blood
35803105|T121|SKI 2053R
35803105|T121|Heptaplatin
35803106|T121|histrelin acetate
35803106|T121|Histrelin
35803107|T121|Hu5F9-G4
35803108|T121|hydrocortisone sodium phosphate
35803108|T121|hydrocortisone sodium succinate
35803108|T121|Hydrocortisone
35803109|T121|dhnp
35803109|T121|hidroxiurea
35803109|T121|hydroxycarbam
35803109|T121|hydroxycarbamid
35803109|T121|hydroxycarbamide
35803109|T121|Hydroxyurea
35803110|T121|IPH 2101
35803111|T121|ibandronate sodium
35803111|T121|ibandronic acid
35803111|T121|Ibandronate
35803112|T121|Ibritumomab tiuxetan
35803113|T121|CRA-032765
35803113|T121|PCI-32765
35803113|T121|Ibrutinib
35803114|T121|BPI-2009H
35803114|T121|Icotinib
35803115|T121|idarubicin comp
35803115|T121|idarubicin hydrochloride
35803115|T121|Idarubicin
35803116|T121|BI 655075
35803116|T121|Idarucizumab
35803117|T121|CAL-101
35803117|T121|GS 1101
35803117|T121|GS-1101
35803117|T121|Idelalisib
35803118|T121|Ifosfamide
35803119|T121|CGP 57148
35803119|T121|CGP57148B
35803119|T121|STI-571
35803119|T121|imatinib mesilate
35803119|T121|imatinib mesylate
35803119|T121|Imatinib
35803120|T121|GRN163L
35803120|T121|Imetelstat
35803121|T121|Indomethacin
35803122|T121|BGJ398
35803122|T121|Infigratinib
35803123|T121|CMC-544
35803123|T121|Inotuzumab ozogamicin
35803124|T121|Interferon alfa-2a
35803125|T121|Interferon alfa-2b
35803126|T121|Interferon gamma-1b
35803127|T121|Iodine-131
35803128|T121|GDC-0068
35803128|T121|RG-7440
35803128|T121|Ipatasertib
35803129|T121|BMS-734016
35803129|T121|MDX-010
35803129|T121|Ipilimumab
35803130|T121|Camptothecin-11
35803130|T121|CPT-11
35803130|T121|U-101440E
35803130|T121|Irinotecan
35803131|T121|MM-398
35803131|T121|MM398
35803131|T121|PEP-02
35803131|T121|PEP02
35803131|T121|Irinotecan liposome
35803132|T121|Iron dextran
35803133|T121|Iron sucrose
35803134|T121|SAR-650984
35803134|T121|isatuximab-irfc
35803134|T121|Isatuximab
35803135|T121|Ro 4-3780
35803135|T121|13-cis-retinoic acid
35803135|T121|13-cis-vitamin A acid
35803135|T121|13-CRA
35803135|T121|cis-retinoic acid
35803135|T121|isotretinoinum
35803135|T121|neovitamin A
35803135|T121|Isotretinoin
35803136|T121|Itraconazole
35803137|T121|AG-120
35803137|T121|Ivosidenib
35803138|T121|BMS-247550
35803138|T121|azaepothilone B
35803138|T121|epothilone B lactam
35803138|T121|Ixabepilone
35803139|T121|MLN2238
35803139|T121|MLN9708
35803139|T121|Ixazomib
35803140|T121|Ketoconazole
35803141|T121|L-glutamine
35803142|T121|Lactulose
35803143|T121|Lamivudine
35803144|T121|lanreotide acetate
35803144|T121|Lanreotide
35803145|T121|Lansoprazole
35803146|T121|GW572016
35803146|T121|Lapatinib
35803147|T121|DN24-02
35803147|T121|Lapuleucel-T
35803148|T121|LOXO-101
35803148|T121|Larotrectinib
35803149|T121|CC-5013
35803149|T121|IMiD-1
35803149|T121|NSC-703813
35803149|T121|Lenalidomide
35803150|T121|Lenograstim
35803151|T121|E7080
35803151|T121|Lenvatinib
35803152|T121|Lepirudin
35803153|T121|CEP-701
35803153|T121|Lestaurtinib
35803154|T121|CGS 20267
35803154|T121|Letrozole
35803155|T121|A-43818
35803155|T121|TAP-144
35803155|T121|leuprolide acetate
35803155|T121|leuprorelin
35803155|T121|leuprorelin acetate
35803155|T121|Leuprolide
35803156|T121|Levamisole
35803157|T121|Levofloxacin
35803158|T121|levoleucovorin calcium
35803158|T121|Levoleucovorin
35803159|T121|XM22
35803159|T121|Lipefilgrastim
35803160|T121|D-19466
35803160|T121|Lobaplatin
35803161|T121|CCNU
35803161|T121|Lomustine
35803162|T121|Loperamide
35803163|T121|Lorazepam
35803164|T121|PF-06463922
35803164|T121|Lorlatinib
35803165|T121|Lusutrombopag
35803166|T121|Lutetium Lu 177 dotatate
35803167|T121|MOR202
35803168|T121|tafasitamab-cxix
35803168|T121|MOR208
35803168|T121|MOR00208
35803168|T121|XmAb5574
35803168|T121|Tafasitamab
35803169|T121|Mannitol
35803170|T121|HGS-ETR1
35803170|T121|Mapatumumab
35803171|T121|AB1010
35803171|T121|Masitinib
35803172|T121|nitrogen mustard
35803172|T121|Mechlorethamine
35803173|T121|medroxyprogesterone acetate
35803173|T121|MPA
35803173|T121|Medroxyprogesterone
35803174|T121|SC10363
35803174|T121|megestrol acetate
35803174|T121|Megestrol
35803175|T121|L-PAM
35803175|T121|L-Sacrolysin
35803175|T121|L-Sarcolysin
35803175|T121|MPL
35803175|T121|phenylalanine mustard
35803175|T121|Melphalan
35803176|T121|Mepolizumab
35803177|T121|6-MP
35803177|T121|6-Mercaptopurine
35803177|T121|Mercaptopurine
35803178|T121|Mesna
35803179|T121|amethopterin
35803179|T121|MTX
35803179|T121|Methotrexate
35803180|T121|8-MOP
35803180|T121|methoxypsoralen
35803180|T121|Methoxsalen
35803181|T121|methylprednisolone acetate
35803181|T121|methylprednisolone sodium succinate
35803181|T121|Methylprednisolone
35803182|T121|Metoclopramide
35803183|T121|PKC412
35803183|T121|Midostaurin
35803184|T121|mitomycin-C
35803184|T121|MTC
35803184|T121|Mitomycin
35803185|T121|o,p′-DDD
35803185|T121|Mitotane
35803186|T121|mitozantrone
35803186|T121|Mitoxantrone
35803187|T121|MGCD0103
35803187|T121|Mocetinostat
35803188|T121|KW-0761
35803188|T121|mogamulizumab-kpkc
35803188|T121|Mogamulizumab
35803189|T121|CYT387
35803189|T121|GS-0387
35803189|T121|Momelotinib
35803190|T121|Montelukast
35803191|T121|AMG 706
35803191|T121|Motesanib
35803192|T121|CAT-8015
35803192|T121|HA22
35803192|T121|moxetumomab pasudotox-tdfk
35803192|T121|Moxetumomab pasudotox
35803193|T121|Mycophenolate mofetil
35803194|T121|NEOD001
35803195|T121|Nabilone
35803196|T121|Nadroparin
35803197|T121|IMC-11F8
35803197|T121|Necitumumab
35803198|T121|254-S
35803198|T121|nedaplat
35803198|T121|Nedaplatin
35803199|T121|506U78
35803199|T121|Nelarabine
35803200|T121|HKI-272
35803200|T121|Neratinib
35803201|T121|NEPA
35803201|T121|Netupitant and palonosetron
35803202|T121|AMN107
35803202|T121|Nilotinib
35803203|T121|Nilutamide
35803204|T121|pimustine
35803204|T121|ACNU
35803204|T121|Nimustine
35803205|T121|BIBF 1120
35803205|T121|Nintedanib
35803206|T121|MK4827
35803206|T121|Niraparib
35803207|T121|MDX-1106
35803207|T121|ONO-4538
35803207|T121|BMS-936558
35803207|T121|Nivolumab
35803208|T121|Nolatrexed
35803209|T121|NPLD
35803209|T121|liposome-encapsulated doxorubicin citrate
35803209|T121|Non-pegylated liposomal doxorubicin
35803210|T121|Norethandrolone
35803211|T121|GA101
35803211|T121|R7159
35803211|T121|RO5072759
35803211|T121|afutuzumab
35803211|T121|Obinutuzumab
35803212|T121|SMS 201-995
35803212|T121|octreotide immediate release
35803212|T121|octreotide IR
35803212|T121|octreotide acetate
35803212|T121|Octreotide
35803213|T121|octreotide acetate for injectable suspension
35803213|T121|octreotide long-acting release
35803213|T121|Octreotide LAR
35803214|T121|HuMax-CD20
35803214|T121|Ofatumumab
35803215|T121|Olanzapine
35803216|T121|AZD-2281
35803216|T121|KU-0059436
35803216|T121|AZD2281
35803216|T121|Olaparib
35803217|T121|LY3012207
35803217|T121|IMC-3G3
35803217|T121|Olaratumab
35803218|T121|homoharringtonine
35803218|T121|omacetaxine mepesuccinate
35803218|T121|HHT
35803218|T121|Omacetaxine
35803219|T121|Omeprazole
35803220|T121|MetMAb
35803220|T121|RO5490258
35803220|T121|Onartuzumab
35803221|T121|SN-307
35803221|T121|Ondansetron
35803222|T121|Oprelvekin
35803223|T121|ONX 0912
35803223|T121|Oprozomib
35803224|T121|TAK-700
35803224|T121|Orteronel
35803225|T121|AZD9291
35803225|T121|Osimertinib
35803226|T121|TRU-016
35803226|T121|Otlertuzumab
35803227|T121|JM-83
35803227|T121|RP-54780
35803227|T121|SR-96669
35803227|T121|Oxaliplatin
35803228|T121|ABI-007
35803228|T121|ab-pac
35803228|T121|ab-paclitaxel
35803228|T121|nab-paclitaxel
35803228|T121|paclitaxel protein-bound
35803228|T121|paclitaxel protein-bound particles for injectable suspension (albumin-bound)
35803228|T121|albumin-bound paclitaxel
35803228|T121|Paclitaxel nanoparticle albumin-bound
35803229|T121|Paclitaxel
35803230|T121|SB1518
35803230|T121|Pacritinib
35803231|T121|PD-0332991
35803231|T121|Palbociclib
35803232|T121|palonosetron HCL
35803232|T121|Palonosetron
35803233|T121|pamidronate disodium omega
35803233|T121|Pamidronate
35803234|T121|ABX-EGF
35803234|T121|clone E7.6.3
35803234|T121|Panitumumab
35803235|T121|panobinostat lactate anhydrous
35803235|T121|LBH589
35803235|T121|Panobinostat
35803236|T121|Pantoprazole
35803237|T121|GW786034B
35803237|T121|Pazopanib
35803238|T121|pegasparaginase
35803238|T121|PEG-L-asparaginase
35803238|T121|peg-asparginase
35803238|T121|Pegaspargase
35803239|T121|Pegfilgrastim-jmdb
35803240|T121|pegylated GCSF
35803240|T121|pegylated granulocyte colony stimulating factor
35803240|T121|pegylated G-CSF
35803240|T121|Pegfilgrastim
35803241|T121|Peginterferon alfa-2a
35803242|T121|PEG-IFN alfa-2b
35803242|T121|pegylated interferon alfa-2b
35803242|T121|SCH 54031
35803242|T121|polyethylene glycol IFN-A2b
35803242|T121|polyethylene glycol interferon alfa-2b
35803242|T121|Peginterferon alfa-2b
35803243|T121|doxorubicin HCl liposome injection
35803243|T121|PLD
35803243|T121|Pegylated liposomal doxorubicin
35803244|T121|lambrolizumab
35803244|T121|MK-3475
35803244|T121|SCH 900475
35803244|T121|Pembrolizumab
35803245|T121|pemetrexed disodium
35803245|T121|Pemetrexed
35803246|T121|pentamidine dimesilate
35803246|T121|Pentamidine
35803247|T121|dCF
35803247|T121|2'-deoxycoformycin
35803247|T121|Pentostatin
35803248|T121|PRM-151
35803248|T121|Pentraxin 2
35803249|T121|KRX-0401
35803249|T121|Perifosine
35803250|T121|Rhumab 2C4
35803250|T121|2C4
35803250|T121|Pertuzumab
35803251|T121|Phenytoin
35803252|T121|vitamin K
35803252|T121|Phytonadione
35803253|T121|GDC-0941
35803253|T121|Pictilisib
35803254|T121|MDV9300
35803254|T121|CT-011
35803254|T121|Pidilizumab
35803255|T121|theprubicin
35803255|T121|1609-RB
35803255|T121|THP-doxorubicin
35803255|T121|Pirarubicin
35803256|T121|BBR 2778
35803256|T121|pixantrone dimaleate
35803256|T121|Pixantrone
35803257|T121|AMD3100
35803257|T121|Plerixafor
35803258|T121|mithramycin
35803258|T121|Plicamycin
35803259|T121|NPI-2358
35803259|T121|Plinabulin
35803260|T121|CC-4047
35803260|T121|3-amino-thalidomide
35803260|T121|CC4047
35803260|T121|Pomalidomide
35803261|T121|ponatinib hydrochloride
35803261|T121|AP24534
35803261|T121|Ponatinib
35803262|T121|Porfimer
35803263|T121|SB939
35803263|T121|Pracinostat
35803264|T121|Pralatrexate
35803265|T121|Prasugrel
35803266|T121|Pravastatin
35803267|T121|delta(1)hydrocortisone
35803267|T121|metacortandralone
35803267|T121|prednisolone acetate
35803267|T121|delta1-dehydro-hydrocortisone
35803267|T121|deltahydrocortisone
35803267|T121|prednisolone tebutate
35803267|T121|Prednisolone
35803268|T121|pred
35803268|T121|Prednisone
35803269|T121|Ro 4-6467/1
35803269|T121|ibenzmethyzine hydrochloride
35803269|T121|NCI-C01810
35803269|T121|procarbazine hydrochloride
35803269|T121|ibenzmethyzin hydrochloride
35803269|T121|P-Carbazine
35803269|T121|Procarbazine
35803270|T121|Prochlorperazine
35803271|T121|Promethazine
35803272|T121|Protamine sulfate
35803273|T121|4-factor prothrombin complex concentrate
35803273|T121|factor IX complex
35803273|T121|PCC
35803273|T121|Prothrombin Complex Concentrate human
35803274|T121|Quinine
35803275|T121|JNJ-26481585
35803275|T121|Quisinostat
35803276|T121|AC220
35803276|T121|ASP2689
35803276|T121|Quizartinib
35803277|T121|Rabeprazole
35803278|T121|Radium Ra 223 dichloride
35803278|T121|Radium-223 chloride
35803278|T121|Ra-223
35803278|T121|Radium-223
35803279|T121|IY5511HCl
35803279|T121|Radotinib
35803280|T121|Raloxifene
35803281|T121|ZD 1694
35803281|T121|raltitrexed disodium
35803281|T121|TDX
35803281|T121|Raltitrexed
35803282|T121|Ramosetron
35803283|T121|LY3009806
35803283|T121|IMC-1121B
35803283|T121|Ramucirumab
35803284|T121|MCNU
35803284|T121|ranomustine
35803284|T121|Ranimustine
35803285|T121|Ranitidine
35803286|T121|Rasburicase
35803287|T121|BAY 869766
35803287|T121|Refametinib
35803288|T121|BAY 73-4506
35803288|T121|Regorafenib
35803289|T121|IPI-504
35803289|T121|Retaspimycin
35803290|T121|Rho(D) immune globulin
35803291|T121|LEE-011
35803291|T121|LEE011
35803291|T121|Ribociclib
35803292|T121|ACY-1215
35803292|T121|rocilinostat
35803292|T121|Ricolinostat
35803293|T121|AMG 102
35803293|T121|Rilotumumab
35803294|T121|Risedronate
35803295|T121|Rituximab-abbs
35803296|T121|IDEC-102
35803296|T121|BI 695500
35803296|T121|RTXM83
35803296|T121|IDEC-C2B8
35803296|T121|PF-05280586
35803296|T121|Rituximab
35803297|T121|Rituximab and hyaluronidase human
35803298|T121|BAY 59-7939
35803298|T121|Rivaroxaban
35803299|T121|CO-1686
35803299|T121|Rociletinib
35803300|T121|SCH-619734
35803300|T121|SCH619734
35803300|T121|Rolapitant
35803301|T121|FR901228
35803301|T121|FK228
35803301|T121|NSC 630176
35803301|T121|depsipeptide
35803301|T121|Romidepsin
35803302|T121|Romiplostim
35803303|T121|AOP2014
35803303|T121|Ropeginterferon alfa-2b
35803304|T121|CO-338
35803304|T121|AG-014699
35803304|T121|PF-0136738
35803304|T121|Rucaparib
35803305|T121|ruxolitinib phosphate
35803305|T121|INCB018424
35803305|T121|Ruxolitinib
35803306|T121|sacituzumab govitecan-hziy
35803306|T121|RS7-SN38
35803306|T121|IMMU-132
35803306|T121|Sacituzumab govitecan
35803307|T121|lexidronam pentasodium
35803307|T121|153-Sm-EDTMP
35803307|T121|153Sm-ethylenediaminetetramethylenephosphonate (EDTMP)
35803307|T121|samarium [153 SM]
35803307|T121|samarium Sm 153 lexidronam injection
35803307|T121|Samarium-153
35803308|T121|CS-682
35803308|T121|Sapacitabine
35803309|T121|GMCSF
35803309|T121|GM-CSF
35803309|T121|granulocyte macrophage colony stimulating factor
35803309|T121|Sargramostim
35803310|T121|Scopolamine
35803311|T121|KPT-330
35803311|T121|Selinexor
35803312|T121|AZD6244
35803312|T121|Selumetinib
35803313|T121|AVE5026
35803313|T121|Semuloparin
35803314|T121|methyl-lomustine
35803314|T121|MeCCNU
35803314|T121|methyl-CCNU
35803314|T121|Semustine
35803315|T121|senna
35803315|T121|Sennosides
35803316|T121|CNTO 328
35803316|T121|Siltuximab
35803317|T121|APC8015
35803317|T121|Sipuleucel-T
35803318|T121|WY-090217
35803318|T121|AY 22989
35803318|T121|SILA 9268A
35803318|T121|rapamycin
35803318|T121|SLM
35803318|T121|RAPA
35803318|T121|Sirolimus
35803319|T121|LDE225
35803319|T121|erismodegib
35803319|T121|Sonidegib
35803320|T121|BAY 54-9085
35803320|T121|BAY 43-9006
35803320|T121|Sorafenib
35803321|T121|CC-292
35803321|T121|AVL-292
35803321|T121|Spebrutinib
35803322|T121|STZ
35803322|T121|Streptozocin
35803323|T121|sunitinib malate
35803323|T121|SU011248
35803323|T121|SU11248
35803323|T121|Sunitinib
35803324|T121|FK-506
35803324|T121|Tacrolimus
35803325|T121|SL-401
35803325|T121|tagraxofusp-erzs
35803325|T121|Tagraxofusp
35803326|T121|BMN-673
35803326|T121|Talazoparib
35803327|T121|T-VEC
35803327|T121|Talimogene laherparepvec
35803328|T121|Tamibarotene
35803329|T121|tamoxifen citrate
35803329|T121|ICI-46474
35803329|T121|TAM
35803329|T121|TMX
35803329|T121|Tamoxifen
35803330|T121|Tbo-filgrastim
35803331|T121|S-1
35803331|T121|Tegafur gimeracil oteracil
35803332|T121|tegafur-uracil
35803332|T121|Tegafur and uracil
35803333|T121|telotristat ethyl as telotristat etiprate
35803333|T121|Telotristat
35803334|T121|TMZ
35803334|T121|Temozolomide
35803335|T121|CCI-779
35803335|T121|Temsirolimus
35803336|T121|VM-26
35803336|T121|Teniposide
35803337|T121|DJ-927
35803337|T121|Tesetaxel
35803338|T121|Thalidomide
35803339|T121|6-thioguanine
35803339|T121|6-TG
35803339|T121|2-Amino-6-Mercaptopurine
35803339|T121|tioguanine
35803339|T121|Thioguanine
35803340|T121|Thiophosphoamide
35803340|T121|TSPA
35803340|T121|TESPA
35803340|T121|Thiotepa
35803341|T121|Ticagrelor
35803342|T121|Ticlopidine
35803343|T121|CS-1008
35803343|T121|Tigatuzumab
35803344|T121|Tinzaparin
35803345|T121|R115777
35803345|T121|Tipifarnib
35803346|T121|Tirofiban
35803347|T121|CTL019
35803347|T121|CART19
35803347|T121|tisagenlecleucel-T
35803347|T121|Tisagenlecleucel
35803348|T121|ARQ 197
35803348|T121|Tivantinib
35803349|T121|AV-951
35803349|T121|Tivozanib
35803350|T121|Tocilizumab
35803351|T121|CP-690550
35803351|T121|tasocitinib
35803351|T121|Tofacitinib
35803352|T121|SKF S-104864-A
35803352|T121|Topotecan
35803353|T121|Toremifene
35803354|T121|CHR-2797
35803354|T121|Tosedostat
35803355|T121|tositumomab and iodine-131 tositumomab
35803355|T121|tositumomab and I 131 tositumomab
35803355|T121|Tositumomab and I-131
35803356|T121|ET-743
35803356|T121|Trabectedin
35803357|T121|GSK-1120212
35803357|T121|GSK1120212
35803357|T121|JTP-74057
35803357|T121|trametinib dimethyl sulfoxide
35803357|T121|Trametinib
35803358|T121|Tranexamic acid
35803359|T121|Trastuzumab-dkst
35803360|T121|CT-P6
35803360|T121|Trastuzumab-pkrb
35803361|T121|Trastuzumab
35803362|T121|AMG 386
35803362|T121|Trebananib
35803363|T121|CP-675
35803363|T121|CP-675206
35803363|T121|ticilimumab
35803363|T121|Tremelimumab
35803364|T121|Treosulfan
35803365|T121|trifluridine/tipiracil
35803365|T121|TAS-102
35803365|T121|trifluridine and tipiracil
35803365|T121|Trifluridine and tipiracil
35803366|T121|co-trimoxazole
35803366|T121|SMZ-TMP
35803366|T121|SMZ-TMP DS
35803366|T121|TMP-SMX
35803366|T121|TMS
35803366|T121|SMX / TMP
35803366|T121|cotrimazole
35803366|T121|cotrimoxazole
35803366|T121|SMZ ( CO )
35803366|T121|Trimethoprim-Sulfamethoxazole
35803367|T121|triptorelin pamoate
35803367|T121|CL118532
35803367|T121|AY25650
35803367|T121|Triptorelin
35803368|T121|ICS 205-930
35803368|T121|Tropisetron
35803369|T121|LFB-R603
35803369|T121|TG-1101
35803369|T121|TGTX-1101
35803369|T121|TG-20
35803369|T121|Ublituximab
35803370|T121|UFH
35803370|T121|Unfractionated heparin
35803371|T121|uramustine
35803371|T121|Uracil mustard
35803372|T121|Uridine triacetate
35803373|T121|33A
35803373|T121|SGN-CD33A
35803373|T121|Vadastuximab talirine
35803374|T121|valaciclovir
35803374|T121|BW-256U
35803374|T121|acyclovir-valine
35803374|T121|valaciclovir Hcl
35803374|T121|ValACV
35803374|T121|Valacyclovir
35803375|T121|Valganciclovir
35803376|T121|valproic acid
35803376|T121|Valproate
35803377|T121|AD 32
35803377|T121|Valrubicin
35803378|T121|AZD6474
35803378|T121|ZD6474
35803378|T121|Vandetanib
35803379|T121|CDX-1127
35803379|T121|Varlilumab
35803380|T121|ABT-888
35803380|T121|Veliparib
35803381|T121|hA20
35803381|T121|IMMU-160
35803381|T121|Veltuzumab
35803382|T121|RO5185426
35803382|T121|PLX4032
35803382|T121|RG7204
35803382|T121|Vemurafenib
35803383|T121|GDC-0199
35803383|T121|ABT-199
35803383|T121|Venetoclax
35803384|T121|vincaleukoblastine
35803384|T121|vinblastine sulfate
35803384|T121|vinblastine sulphate
35803384|T121|VLB
35803384|T121|chlorhexamide
35803384|T121|Vinblastine
35803385|T121|VCR
35803385|T121|leurocristine
35803385|T121|vincristine sulfate
35803385|T121|LCR
35803385|T121|Vincristine
35803386|T121|VSLI
35803386|T121|vincristine sulfate liposome injection
35803386|T121|Vincristine liposomal
35803387|T121|LY-099094
35803387|T121|desacetylvinblastine amide
35803387|T121|DVA
35803387|T121|VDS
35803387|T121|DAVA
35803387|T121|Vindesine
35803388|T121|Vinflunine
35803389|T121|KW-2307
35803389|T121|NVB
35803389|T121|vinorelbine tartrate
35803389|T121|Vinorelbine
35803390|T121|GDC-0449
35803390|T121|Vismodegib
35803391|T121|BI 6727
35803391|T121|Volasertib
35803392|T121|Vorapaxar
35803393|T121|Voriconazole
35803394|T121|Vorinostat
35803395|T121|voreloxin
35803395|T121|SNS-595
35803395|T121|Vosaroxin
35803396|T121|warfarina sodica
35803396|T121|Warfarin
35803397|T121|azidothymidine
35803397|T121|AZT
35803397|T121|ZDV
35803397|T121|Zidovudine
35803398|T121|VEGF trap
35803398|T121|aflibercept
35803398|T121|Ziv-aflibercept
35803399|T121|acido zoledronico
35803399|T121|zoledronate
35803399|T121|Zoledronic acid
42542125|T121|Acquired coagulopathy
42542126|T121|Acute myeloid leukemia
42542127|T121|Acute promyelocytic leukemia
42542128|T121|Carcinoma of unknown primary
42542129|T121|Adrenocortical carcinoma
42542130|T121|Adult T-cell leukemia-lymphoma
42542131|T121|Allogeneic HSCT
42542132|T121|Anal cancer
42542133|T121|Anaplastic glioma
42542134|T121|Anaplastic large cell lymphoma
42542135|T121|Antiphospholipid antibody syndrome
42542136|T121|Aplastic anemia
42542137|T121|Atypical hemolytic uremic syndrome
42542138|T121|Autoimmune cytopenia
42542139|T121|Warm autoimmune hemolytic anemia
42542140|T121|Autologous HSCT
42542141|T121|B-cell acute lymphoblastic leukemia
42542142|T121|Bladder cancer
42542143|T121|Blastic plasmacytoid dendritic cell neoplasm
42542144|T121|Bone sarcoma
42542145|T121|Breast cancer
42542146|T121|Burkitt lymphoma
42542147|T121|CNS carcinoma
42542148|T121|CNS leukemia
42542149|T121|CNS lymphoma
42542150|T121|CNS melanoma
42542151|T121|Castleman disease
42542152|T121|Cervical cancer
42542153|T121|Cholangiocarcinoma
42542154|T121|Chronic lymphocytic leukemia
42542155|T121|Chronic myeloid leukemia
42542156|T121|Chronic myelomonocytic leukemia
42542157|T121|Cold agglutinin disease
42542158|T121|Colon cancer
42542159|T121|Cutaneous T-cell lymphoma
42542160|T121|Cutaneous basal cell carcinoma
42542161|T121|Cutaneous squamous cell carcinoma
42542162|T121|Diffuse large B-cell lymphoma
42542163|T121|Endometrial cancer
42542164|T121|Erdheim-Chester disease
42542165|T121|Esophageal cancer
42542166|T121|Essential thrombocythemia
42542167|T121|Ewing sarcoma
42542168|T121|Extranodal NK- and T-cell lymphoma nasal type
42542169|T121|Follicular lymphoma
42542170|T121|Gallbladder cancer
42542171|T121|Gastric cancer
42542172|T121|Gastrointestinal stromal tumor
42542173|T121|Gestational trophoblastic neoplasia
42542174|T121|Glioblastoma
42542175|T121|Graft versus host disease
42542176|T121|HIV-associated lymphoma
42542177|T121|Hairy cell leukemia
42542178|T121|Head and neck cancer
42542179|T121|Hemophagocytic lymphohistiocytosis
42542180|T121|Heparin-induced thrombocytopenia
42542181|T121|Hepatoblastoma
42542182|T121|Hepatocellular carcinoma
42542183|T121|Hereditary hemorrhagic telangiectasia
42542184|T121|Hodgkin lymphoma
42542185|T121|Hodgkin lymphoma nodular lymphocyte-predominant
42542186|T121|Hypereosinophilic syndrome
42542187|T121|Immune thrombocytopenia
42542188|T121|Inherited coagulopathy
42542189|T121|Inherited thrombophilia
42542190|T121|Langerhans cell histiocytosis
42542191|T121|Large granular lymphocytic leukemia
42542192|T121|Light-chain (AL) amyloidosis
42542193|T121|Low-grade glioma
42542194|T121|Mismatch repair deficient malignancy
42542195|T121|Mantle cell lymphoma
42542196|T121|Marginal zone lymphoma
42542197|T121|Mediastinal gray-zone lymphoma
42542198|T121|Medulloblastoma
42542199|T121|Melanoma
42542200|T121|Meningioma
42542201|T121|Merkel cell carcinoma
42542202|T121|Mesothelioma
42542203|T121|Multiple myeloma
42542204|T121|Myelodysplastic syndrome
42542205|T121|Myelofibrosis
42542206|T121|NET of unknown primary
42542207|T121|NK- and T-cell lymphoma
42542208|T121|Nasopharyngeal carcinoma
42542209|T121|Neuroblastoma
42542210|T121|Neuroendocrine tumor
42542211|T121|Non-small cell lung cancer
42542212|T121|Oropharyngeal cancer
42542213|T121|Osteosarcoma
42542214|T121|Ovarian cancer
42542215|T121|POEMS syndrome
42542216|T121|Pancreatic NET
42542217|T121|Pancreatic cancer
42542218|T121|Paroxysmal nocturnal hemoglobinuria
42542219|T121|Penile cancer
42542220|T121|Periampullary adenocarcinoma
42542221|T121|Peripheral T-cell lymphoma
42542222|T121|Pheochromocytoma
42542223|T121|Plasma cell leukemia
42542224|T121|Polycythemia vera
42542225|T121|Post-transplant lymphoproliferative disorder
42542226|T121|Primary mediastinal B-cell lymphoma
42542227|T121|Prostate cancer
42542228|T121|Rectal cancer
42542229|T121|Renal cell carcinoma
42542230|T121|Rhabdomyosarcoma
42542231|T121|Rosai-Dorfman-Destombes disease
42542232|T121|SCC of unknown primary
42542233|T121|Sickle cell anemia
42542234|T121|Small cell lung cancer
42542235|T121|Soft tissue sarcoma
42542236|T121|Stem cell mobilization
42542237|T121|Systemic mastocytosis
42542238|T121|T-cell acute lymphoblastic leukemia
42542239|T121|Testicular cancer
42542240|T121|Thrombocytopenia in liver disease
42542241|T121|Thrombotic thrombocytopenic purpura
42542242|T121|Thymoma
42542243|T121|Thyroid cancer
42542244|T121|Transformed lymphoma
42542245|T121|Uveal melanoma
42542246|T121|Vascular sarcoma
42542247|T121|Venous thromboembolism
42542248|T121|Vulvar cancer
42542249|T121|WHIM syndrome
42542250|T121|Waldenstroem macroglobulinemia
42542251|T121|Wilms tumor
35803400|T121|Anticoagulation
35803401|T121|Chemotherapy
35803402|T121|Chemohormonotherapy
35803403|T121|Chemoimmunotherapy
35803404|T121|Chemoradiotherapy
35803405|T121|Chemoradioimmunotherapy
35803406|T121|Growth factor therapy
35803407|T121|Endocrine therapy
35803408|T121|Hormonoradiotherapy
35803409|T121|Immunosuppressive therapy
35803410|T121|Immunotherapy
35803411|T121|Radiotherapy
35803412|T121|Radioconjugate therapy
35803413|T121|Supportive therapy
35803414|T121|Clotinab
35803415|T121|ReoPro
35803416|T121|Verzenio
35803417|T121|Zytiga
35803418|T121|Calquence
35803419|T121|Calpol
35803420|T121|Panadol
35803421|T121|Tylenol
35803422|T121|Aclacin
35803423|T121|Aclacinomycine
35803424|T121|Aclacinon
35803425|T121|Aclaplastin
35803426|T121|Jaclacin
35803427|T121|All lines of therapy
35803428|T121|Cyclophosphamide and Prednisolone
35803429|T121|Cyclophosphamide and Prednisone
35803429|T121|CP
35803429|T121|CyPred
35803430|T121|Prednisone monotherapy
35803431|T121|Prednisolone monotherapy
35803432|T121|Rituximab monotherapy
35803433|T121|Induction therapy
35803434|T121|7 plus 3d
35803435|T121|High-dose Cytarabine monotherapy (HiDAC)
35803435|T121|HiDAC
35803435|T121|High Dose Ara-C (Cytarabine)
35803435|T121|HDAC
35803435|T121|HDAraC
35803435|T121|High Dose AraC (Cytarabine)
35803436|T121|Intermediate-dose Cytarabine monotherapy (IDAC)
35803436|T121|IDAC
35803436|T121|Intermediate Dose Ara-C (Cytarabine)
35803436|T121|mIDAC
35803436|T121|modified Intermediate Dose Ara-C (Cytarabine)
911923|T121|Aminoblastin
911924|T121|Antiestrogen
911925|T121|Capecitabine and Trastuzumab (XH) and Tucatinib
35803437|T121|7 plus 3d (intermediate-dose)
35803437|T121|7 days of cytarabine + 3 days of daunorubicin
35803438|T121|Granulocyte colony-stimulating factors
35803439|T121|5 plus 2d
35803440|T121|CLAG
35803440|T121|CLadribine, Ara-C (Cytarabine), G-CSF
35803441|T121|HAM
35803441|T121|High-dose Ara-C (Cytarabine), Mitoxantrone
35803441|T121|NOAC
35803441|T121|High-dose Ara-C (Cytarabine) and Mitoxantrone
35803441|T121|NOvantrone (Mitoxantrone) and Ara-C (Cytarabine)
35803442|T121|Cytarabine and Daunorubicin
911926|T121|CapeOx and Erlotinib
911926|T121|Capecitabine, OXaliplatin, Erlotinib
35102032|T121|AspaMetDex (Erwinaze)
35102032|T121|Asparaginase, Methotrexate, Dexamethasone
911927|T121|Contergan
35803444|T121|7 plus 3d (high-dose)
35803444|T121|7 days of cytarabine + 3 days of daunorubicin
35803445|T121|7 plus 3d and GO
35803445|T121|7+3d and GO
35803445|T121|7 days of Cytarabine, 3 days of daunorubicin, Gemtuzumab Ozogamicin
35803446|T121|Cytarabine, Daunorubicin, Gemtuzumab ozogamicin
35803447|T121|7 plus 3i
35803447|T121|7+3i
35803447|T121|7 days of cytarabine + 3 days of idarubicin
35803447|T121|AI
35803447|T121|IA
35803447|T121|Ara-C (Cytarabine) and Idarubicin
35803447|T121|Idarubicin and Ara-C (Cytarabine)
35803443|T121|Cytarabine and Idarubicin
35803448|T121|CYVE
35803448|T121|CYtarabine and VEpesid (Etoposide)
35803448|T121|CYtarabine and VEpeside (Etoposide)
35803448|T121|CYtarabine, VEpesid (Etoposide)
35803448|T121|EA
35803448|T121|Etoposide and Ara-C (Cytarabine)
35102031|T121|BEACOPP-14 (Prednisolone)
35102031|T121|Bleomycin, Etoposide, Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Procarbazine, Prednisolone, 14-day course
911928|T121|Detryptoreline
911929|T121|Distaval
911930|T121|Drugs by local effect
911931|T121|Elipten
35803449|T121|7 plus 3i and Sorafenib
35803450|T121|Cytarabine, Idarubicin, Sorafenib
35803451|T121|7 plus 3d and Glasdegib
35803452|T121|7 plus 3m
35803452|T121|7+3m
35803452|T121|7 days of cytarabine + 3 days of mitoxantrone
35803452|T121|Mitoxantrone and Ara-C (Cytarabine)
35803453|T121|ADE (standard-dose Ara-C)
35803453|T121|ADE
35803453|T121|7-3-7
35803453|T121|8-3-5
35803453|T121|10-3-5
35803453|T121|Ara-C (Cytarabine), Daunorubicin, Etoposide
35803453|T121|7 days of Cytarabine, 3 days of Daunorubicin, 7 days of Etoposide
35803453|T121|8 days of Cytarabine, 3 days of Daunorubicin, 5 days of Etoposide
35803453|T121|10 days of Cytarabine, 3 days of Daunorubicin, 5 days of Etoposide
911932|T121|Farestone
35803454|T121|ADE (high-dose Ara-C)
35803454|T121|ADE
35803454|T121|HIDAC-3-5
35803454|T121|HIDAC-3-7
35803454|T121|Ara-C (Cytarabine), Daunorubicin, Etoposide
35803454|T121|HIgh-Dose Ara-C (Cytarabine), 3 days of Daunorubicin, 5 days of Etoposide
35803454|T121|HIgh-Dose Ara-C (Cytarabine), 3 days of Daunorubicin, 7 days of Etoposide
35803455|T121|CIA
35803455|T121|Clofarabine, Idarubicin, Ara-C (Cytarabine)
35807523|T121|DA 3  plus  10, GO
35807523|T121|DA 3 + 10, GO
35807523|T121|Daunorubicin and Ara-C (Cytarabine), 3 days of daunorubicin + 10 days of cytarabine, Gemtuzumab Ozogamicin
35807524|T121|DA 3  plus  10
35807524|T121|DA 3 + 10
35807524|T121|Da unorubicin and Ara-C (Cytarabine), 3 days of daunorubicin + 10 days of cytarabine
35807524|T121|Daunorubicin and Ara-C (Cytarabine), 3 days of daunorubicin + 10 days of cytarabine
35102030|T121|Carboplatin and Cisplatin
35102030|T121|CC
35102030|T121|Cisplatin and Carboplatin
35803456|T121|DAC
35803456|T121|Daunorubicin, Ara-C (Cytarabine), Cladribine
35803457|T121|FLAG-Ida
35803457|T121|FLudarabine, Ara-C (Cytarabine), G-CSF (Filgrastim), Idarubicin
35803457|T121|FLudarabine, Ara-C (Cytarabine), G-CSF (Lenograstim), Idarubicin
35803458|T121|HAA
35803458|T121|Homoharringtonine (Omacetaxine), Ara-C (Cytarabine), Aclarubicin
35803459|T121|HAD
35803459|T121|Homoharringtonine (Omacetaxine), Ara-C (Cytarabine), Daunorubicin
35803460|T121|AIE
35803460|T121|Ara-C (Cytarabine), Idarubicin, Etoposide
35803460|T121|Idarubicin, Cytarabine, Etoposide
42542252|T121|Adakveo
911933|T121|FUOX and RT
911933|T121|FluoroUracil, OXaliplatin, Radiation Therapy
35803461|T121|ICL
35803461|T121|Idarubicin, Cytarabine, Lomustine
35803462|T121|IC and Norethandrolone/6-MP, MTX, Norethandrolone
35803462|T121|Idarubicin, Cytarabine, Norethandrolone
35803463|T121|MEC
35803463|T121|Mitoxantrone, Etoposide, Cytarabine
35803463|T121|MICE
35803463|T121|MAE
35803463|T121|MItoxantrone, Cytarabine, Etoposide
35803463|T121|Mitoxantrone, Ara-C (Cytarabine), Etoposide
42542253|T121|Anti-nectin-4 antibody
911934|T121|Acalabrutinib and Obinutuzumab
35803464|T121|Non-curative first-line induction therapy
35803465|T121|Azacitidine monotherapy
35803466|T121|Azacitidine and Venetoclax
35803467|T121|Azacitidine and Gemtuzumab ozogamicin
35803468|T121|Best supportive care
35102029|T121|CEOP (Prednisolone)
35102029|T121|Cyclophosphamide, Epirubicin, Oncovin (Vincristine), Prednisolone
35102028|T121|CHOP (Prednisolone)
35102028|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisolone
35803469|T121|Clofarabine monotherapy
35102027|T121|CHOP Modified (Prednisolone)
35102027|T121|mCHOP
35102027|T121|modified Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisolone
35803470|T121|Clofarabine and LoDAC
35803470|T121|Clofarabine and Low Dose Ara-C (Cytarabine)
35803471|T121|Decitabine monotherapy
35803472|T121|Clofarabine and LoDAC/Decitabine
35803472|T121|Clofarabine and Low Dose Ara-C (Cytarabine) alternating with Decitabine
35803473|T121|CPX-351 monotherapy
35803473|T121|Liposomal Cytarabine and Daunorubicin
35102026|T121|CNOP (Prednisolone)
35102026|T121|MCOP
35102026|T121|Cyclophosphamide, Novantrone (Mitoxantrone), Oncovin (Vincristine), Prednisolone
35102026|T121|Mitoxantrone, Cyclophosphamide, Oncovin (Vincristine), Prednisolone
35803474|T121|Decitabine and Venetoclax
35803475|T121|Gemtuzumab ozogamicin monotherapy
35803476|T121|Glasdegib and LoDAC
35803476|T121|Glasdegib and Low Dose Ara-C (Cytarabine)
35803477|T121|Low-dose Cytarabine monotherapy (LoDAC)
35803477|T121|LoDAC
35803477|T121|LDAC
35803477|T121|Low Dose Ara-C (cytarabine)
35803477|T121|Low Dose Ara-C (Cytarabine)
35803477|T121|Low-dose Ara-C (Cytarabine)
35803478|T121|LoDAC and Venetoclax
35803478|T121|Low Dose Ara-C (Cytarabine) and Venetoclax
35803479|T121|Temozolomide monotherapy
35803480|T121|Consolidation after upfront therapy
35803481|T121|Cytarabine and Mitoxantrone (MC)
35803481|T121|MC
35803481|T121|Mitoxantrone and Cytarabine
35803482|T121|Observation
35102025|T121|CVP (Prednisolone)
35102025|T121|Cyclophosphamide, Oncovin (Vincristine), Prednisolone
35803483|T121|HiDAC and G-CSF
35803483|T121|High Dose Ara-C (Cytarabine) and Granulocyte Colony Stimulating Factor
35803484|T121|BuCy
35102024|T121|CVP (Vinblastine/Prednisolone)
35102024|T121|Cyclophosphamide, Vinblastine, Prednisolone
35803485|T121|BuFlu, then allo HSCT
35803485|T121|BuFlu
35803485|T121|Flu/Bu
35803485|T121|Fludarabine and Busulfan
35102023|T121|Cyclophosphamide, Daunorubicin, Vincristine, Prednisolone
35803486|T121|CLARA
35803486|T121|CLofarabine and ARA-C (Cytarabine)
35803486|T121|GCLAC
35803486|T121|G-CSF, Clofarabine, Ara-C (Cytarabine)
35803487|T121|Sorafenib monotherapy
35803488|T121|Cyclophosphamide and TBI, then allo HSCT
35803488|T121|Cy/TBI
35803488|T121|Cyclophosphamide and Total Body Irradiation
35803489|T121|External beam radiotherapy
35803490|T121|Etoposide and Mitoxantrone
35803490|T121|Mitoxantrone and Etoposide
35803491|T121|Fludarabine and TBI, then allo HSCT
35803492|T121|Cyclosporines
35803493|T121|Fludarabine, Busulfan, ATG, then allo HSCT
35803494|T121|CLAG-M
35803494|T121|CLadribine, Ara-C (Cytarabine), G-CSF, Mitoxantrone
35803495|T121|Low-dose TBI, then allo HSCT
35803495|T121|Total Body Irradiation
35803496|T121|Non-curative first-line maintenance therapy
35803497|T121|Salvage therapy
35803498|T121|Clofarabine and Cytarabine
35803499|T121|Serotonin 5-HT3 antagonists
35803500|T121|Clofarabine and Melphalan, then allo HSCT
35102022|T121|Docetaxel and Prednisolone
35102021|T121|DOLP (Prednisolone)
35102021|T121|Daunorubicin, Oncovin (Vincristine), L-Asparaginase, Prednisolone
35102020|T121|eBEACOPP (Prednisolone)
35102020|T121|escalated Bleomycin, Etoposide, Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Procarbazine, Prednisolone
35803501|T121|FLAG
35803501|T121|FLudarabine, Ara-C (Cytarabine), G-CSF
35803502|T121|Cytarabine and Thioguanine
35803503|T121|F-SHAI
35803503|T121|Fludarabine, Sequential High-dose Ara-C (cytarabine), Idarubicin
42542254|T121|Brukinsa
35803504|T121|Consolidation after salvage therapy
35803505|T121|BuCy, then allo HSCT
35803506|T121|FLAG-DNX
35803506|T121|FLudarabine, Ara-C (Cytarabine), G-CSF, DauNoXome (Daunorubicin liposomal)
35803507|T121|Non-curative subsequent-line therapy
35803508|T121|Ruxolitinib monotherapy
35803509|T121|7 plus 3d and Midostaurin
35803509|T121|7+3d and Midostaurin
35803509|T121|7 days of cytarabine, 3 days of daunorubicin, Midostaurin
35803510|T121|HiDAC and Midostaurin
35803510|T121|High Dose Ara-C (Cytarabine) and Midostaurin
42542255|T121|FLT3-positive Acute myeloid leukemia
35803511|T121|7 plus 3d and Sorafenib
35803512|T121|IDAC and Sorafenib
35803512|T121|Intermediate Dose Ara-C (Cytarabine) and Sorafenib
35803513|T121|Midostaurin monotherapy
35803514|T121|Maintenance after upfront therapy
35803515|T121|Gilteritinib monotherapy
35803516|T121|Azacitidine and Sorafenib
35803517|T121|Ivosidenib monotherapy
42542256|T121|IDH-mutated Acute myeloid leukemia
35803518|T121|Enasidenib monotherapy
35803519|T121|5 plus 3d
35803519|T121|5+3d
35803519|T121|5 days of cytarabine + 3 days of daunorubicin
35803520|T121|5 plus 3i
35803520|T121|5+3i
35803520|T121|5 days of cytarabine + 3 days of idarubicin
35803521|T121|7 plus 3d (low-dose)
35803521|T121|7 days of cytarabine + 3 days of daunorubicin
35803522|T121|7 plus 3i and Panobinostat
35803522|T121|7+3i and Panobinostat
35803522|T121|7 days of cytarabine + 3 days of idarubicin, Panobinostat
35803523|T121|Panobinostat monotherapy
35803524|T121|7 plus 3i and Vorinostat
35803525|T121|Cytarabine, Idarubicin, Vorinostat
35803526|T121|7 plus 5i
35803526|T121|7+5i
35803526|T121|7 days of cytarabine + 5 days of idarubicin
35803527|T121|Cytarabine, Daunorubicin, Vincristine
35803528|T121|Cytarabine, Daunorubicin, Mercaptopurine, Prednisolone
35803529|T121|Cytarabine, Doxorubicin, Vincristine, Prednisolone
35803530|T121|Daunorubicin monotherapy
35803531|T121|DAT
35803531|T121|TAD9
35803531|T121|Daunorubicin, Ara-C (Cytarabine), Thioguanine
35803531|T121|Thioguanine, Ara-C (Cytarabine), Daunorubicin
35803531|T121|Thioguanine, Ara-C (Cytarabine), Daunorubicin over 9 days
35102019|T121|FULV/FULV and RT
35102019|T121|FluoroUracil and LeucoVorin (Folinic acid) alternating with FluoroUracil, LeucoVorin (Folinic acid) and Radiation Therapy
35803532|T121|DCTER
35803532|T121|Dexamethasone, Cytarabine, Thioguanine, Etoposide, Rubidomycin (Daunomycin)
35803533|T121|D-ZAPO
35803533|T121|Daunomycin, 5-Azacytidine, Ara-C (Cytarabine), Prednisone, Oncovin (Vincristine)
35803534|T121|Decitabine and Valproate
35803535|T121|Mercaptopurine monotherapy
35803536|T121|PATCO
35803536|T121|Prednisone, Ara-C (Cytarabine), Thioguanine, Cyclophosphamide, Oncovin (Vincristine)
35803537|T121|VAMP (Amethopterin)
35803537|T121|Vincristine, Amethopterin (Methotrexate), Mercaptopurine, Prednisone
35803538|T121|Amsacrine and Cytarabine
35803539|T121|Cytarabine monotherapy
35803540|T121|Vorinostat monotherapy
35803541|T121|POMP
35803541|T121|Purinethol (Mercaptopurine), Oncovin (Vincristine), Methotrexate, Prednisone
35803542|T121|IAP
35803542|T121|Idarubicin, Ara-C (cytarabine), Pravastatin
35803543|T121|SHAI
35803543|T121|Sequential High-dose Ara-C (Cytarabine), Idarubicin
35803544|T121|Vosaroxin and Cytarabine
35803545|T121|Azacitidine, Vorinostat, Gemtuzumab ozogamicin
35803546|T121|Cladribine monotherapy
35803547|T121|ADE and ATRA
35803547|T121|Ara-C (Cytarabine), Daunorubicin, Etoposide, All-Trans Retinoic Acid
35803548|T121|Arsenic trioxide monotherapy
35803549|T121|Arsenic trioxide and ATRA
35803550|T121|Arsenic trioxide, ATRA, Gemtuzumab ozogamicin
35803551|T121|Arsenic trioxide, ATRA, Idarubicin
35803552|T121|ATRA monotherapy
35803553|T121|ATRA, Cytarabine, Daunorubicin
35803554|T121|Arsenic trioxide, then ATRA and Daunorubicin
35803555|T121|ATRA and Daunorubicin
35803556|T121|ATRA, Cytarabine, Idarubicin
35803557|T121|ATRA and Idarubicin
35803557|T121|AIDA
35803557|T121|ATRA, IDArubicin
35803558|T121|Idarubicin, then Mitoxantrone, then Idarubicin
35803559|T121|Cytarabine and Idarubicin, then Etoposide and Mitoxantrone, then Cytarabine, Idarubicin, Thioguanine
35803560|T121|Idarubicin, then Mitoxantrone, then Idarubicin, with ATRA
35803562|T121|Cytarabine and Idarubicin, then Mitoxantrone, then Cytarabine and Idarubicin, with ATRA
35803563|T121|Cytarabine and Idarubicin, then Etoposide and Mitoxantrone, then Cytarabine, Idarubicin, Thioguanine, with ATRA
35803564|T121|ATRA, Mercaptopurine, Methotrexate
35803565|T121|Mercaptopurine and Methotrexate
35803566|T121|Arsenic trioxide and Idarubicin
35803567|T121|Tamibarotene monotherapy
35803568|T121|Cytarabine and G-CSF
35803569|T121|Busulfan and Melphalan, then auto HSCT
35803570|T121|BEP
35803570|T121|PEB
35803570|T121|Bleomycin, Etoposide, Platinol (Cisplatin)
35803570|T121|Platinol (Cisplatin), Etoposide, Bleomycin
35803570|T121|PVP16B
35803570|T121|Platinol (Cisplatin), VP-16 (Etoposide), Bleomycin
35803571|T121|Carboplatin and Docetaxel
35803571|T121|CbD
35803571|T121|DCb
35803571|T121|Docetaxel and Carboplatin
35803572|T121|Carboplatin and Paclitaxel (CP)
35803572|T121|PCb
35803572|T121|Paclitaxel and Carboplatin
35803572|T121|TC
35803572|T121|Taxol (Paclitaxel) and Carboplatin
35803572|T121|CP
35803572|T121|PC
35803572|T121|Carboplatin and Paclitaxel
35803573|T121|Cisplatin monotherapy
35803574|T121|Cisplatin and Docetaxel (DC)
35803574|T121|Taxotere (Docetaxel) and Platinol (Cisplatin)
35803574|T121|TC
35803574|T121|Docetaxel, Cisplatin
35803574|T121|Taxotere (Docetaxel), Cisplatin
35803574|T121|DP
35803574|T121|Doc-Cis
35803574|T121|Docetaxel and Cisplatin
35803574|T121|Docetaxel and Platinol (Cisplatin)
35803574|T121|CD
35803574|T121|Cisplatin and Docetaxel
35803575|T121|Cisplatin and Gemcitabine (GC)
35803575|T121|GC
35803575|T121|Gemcitabine, Cisplatin
35803575|T121|GP
35803575|T121|"<table class=""wikitable"" style=""color:white; background-color:#9e4244"">"
35803575|T121|Gemcitabine and Cisplatin
35803575|T121|Gemcitabine and Platinol (Cisplatin)
35803576|T121|Cisplatin and Irinotecan (IC)
35803576|T121|IC
35803576|T121|Irinotecan and Cisplatin
35803576|T121|CI
35803576|T121|Irinotecan and Platinol (Cisplatin)
35803576|T121|Irinotecan, Platinol (Cisplatin)
35803577|T121|Docetaxel and Gemcitabine
35803577|T121|GD
35803577|T121|GDoc
35803577|T121|Gemcitabine and Docetaxel
35803577|T121|DG
35803578|T121|Steroids
35803579|T121|Erlotinib and Bevacizumab
35803580|T121|GCP
35803580|T121|Gemcitabine, Carboplatin, Paclitaxel
35803580|T121|Gefitinib, Carboplatin, Pemetrexed
35803581|T121|Gemcitabine and Irinotecan
35803582|T121|PCE
35803582|T121|Paclitaxel, Carboplatin, Etoposide
35803582|T121|Taxol (Paclitaxel) Etoposide), Carboplatin
35803583|T121|Kadcyla
35803584|T121|Adjuvant therapy
35803585|T121|Mitotane monotherapy
35803586|T121|Adrenalectomy
35803587|T121|Mitotane and Streptozocin
35803588|T121|Non-curative therapy
35803589|T121|Mitotane and EDP
35803589|T121|Mitotane, Etoposide, Doxorubicin, Platinol (Cisplatin)
35803590|T121|Placebo
35803591|T121|CHOP-14
35803591|T121|CHOP-DI
35803591|T121|I-CHOP
35803591|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne every 14 days
35803591|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne, Dose-Intense
35803591|T121|Intensive Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
35803591|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone, Dose Intense
35803591|T121|Intensified Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone
35803591|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone every 14 days
35803592|T121|Interferon alfa-2b and Zidovudine
35803593|T121|LSG15
35803594|T121|mLSG15
35803595|T121|Alemtuzumab monotherapy
35803596|T121|Lenalidomide monotherapy
35803597|T121|Afanix
35803598|T121|Gilotrif
35803599|T121|Giotrif
35803600|T121|Tomtovok
35803601|T121|Tovok
35803602|T121|Xovoltib
35803603|T121|Macrolin
35803604|T121|Proleukin
35803605|T121|Alecensa
35803606|T121|Campath
35803607|T121|Campath-1H
35803608|T121|Lemtrada
35803609|T121|Mabcampath
35803610|T121|BuCyTBI
35803610|T121|Busulfan, Cyclophosphamide, Total Body Irradiation
35803611|T121|Busulfan and Cyclophosphamide
35803612|T121|Busulfan and Fludarabine
35803612|T121|BuFlu
35803612|T121|Flu/Bu
35803612|T121|Fludarabine and Busulfan
35803613|T121|Cyclophosphamide and TBI
35803613|T121|Cy/TBI
35803613|T121|Cyclophosphamide and Total Body Irradiation
35803613|T121|CY/TBI
35803613|T121|CYclophosphamide and Total Body Irradiation
35102018|T121|Jiebaishu
35803614|T121|Etoposide and TBI
35803614|T121|Etoposide and Total Body Irradiation
35803615|T121|Fludarabine, Busulfan, Cyclophosphamide
35803615|T121|FluBuCy
35803616|T121|BEAM
35803616|T121|BCNU (Carmustine), Etoposide, Ara-C (Cytarabine), Melphalan
35803616|T121|BiCNU (Carmustine), Etoposide, Ara-C (Cytarabine), Melphalan
35803616|T121|Rituximab, BiCNU (Carmustine), Etoposide, Ara-C (Cytarabine), Melphalan
911935|T121|Abiraterone and Enzalutamide
35803617|T121|BFR
35803617|T121|Bendamustine, Fludarabine, Rituximab
35803618|T121|Clofarabine and Melphalan
35803619|T121|Cyclophosphamide, Fludarabine, Thiotepa
35803620|T121|FC
35803620|T121|Fludarabine and Cyclophosphamide
35803620|T121|Fludarabine, Cyclophosphamide
35803620|T121|CF
35803620|T121|Cyclophosphamide and Fludarabine
35803621|T121|FCR
35803621|T121|Fludarabine, Cyclophosphamide, Rituximab
35803621|T121|R-FC
35803621|T121|Rituximab, Fludarabine, Cyclophosphamide
35803621|T121| R-FC
35102017|T121|MCP (Prednisolone)
35102017|T121|Mitoxantrone, Chlorambucil, Prednisolone
35803622|T121|Fludarabine and TBI
911936|T121|AC and Pembrolizumab
911936|T121|Adriamycin (Doxorubicin), Cyclophosphamide, Pembrolizumab
35102016|T121|Mitoxantrone, Asparaginase Erwinia chrysanthemi, Vincristine, Dexamethasone
35803623|T121|Fludarabine, Busulfan, ATG
35803624|T121|Antithymocyte globulin
35102015|T121|MP (Prednisolone)
35102015|T121|MP
35102015|T121|Melphalan and Prednisolone
35803625|T121|Fludarabine, Busulfan, ATG, Ibritumomab tiuxetan
35803626|T121|Fludarabine, Cyclophosphamide, ATG
35803627|T121|Fludarabine, Cyclophosphamide, TBI for dUCB or haploidentical transplant
35803627|T121|dUCB
35803627|T121|double Umbilical Cord Blood
35803628|T121|Fludarabine and Melphalan
35803628|T121|Flu-Mel
35803629|T121|Fludarabine, Melphalan, Alemtuzumab
35803630|T121|Low-dose TBI
35803630|T121|Total Body Irradiation
35803631|T121|TLI and ATG
35803631|T121|Total Lymphocyte Irradiation and Anti-Thymocyte Globulin
35803632|T121|(90)YFC
35803632|T121|Ibritumomab tiuxetan, Fludarabine, Cyclophosphamide
35803633|T121|Abloric
35803634|T121|Aloprim
35803635|T121|Caplenal
35803636|T121|Milurit
35803637|T121|Zyloprim
35803638|T121|Zyloric
35803639|T121|Zyoway
35803640|T121|Actazolam
35803641|T121|Alam-PH
35803642|T121|Alcalm
35803643|T121|Alplax
35803644|T121|Apazol
35803645|T121|Azom
35803646|T121|Azor
35803647|T121|Copax
35803561|T121|Frixitas
35803648|T121|Onax
35803649|T121|Pinix
35803650|T121|Tafil
35803651|T121|Tranax
35803652|T121|Xanax
35803653|T121|Xanor
35803654|T121|Hexalen
35803655|T121|Hexastat
35803656|T121|Cytofos
35803657|T121|Ethyol
35803658|T121|Amicar
35803659|T121|Cytadren
35803660|T121|Orimeten
35803661|T121|Orimetene
35803662|T121|Calsed
35803663|T121|Amekrin
35803664|T121|Amsa P-D
35803665|T121|Amsidine
35803666|T121|Amsidyl
35803667|T121|Lamasine
35803668|T121|Agrylin
35803669|T121|Xagrid
35803670|T121|Definitive therapy
35803671|T121|Capecitabine, Mitomycin, RT
911937|T121|ADE and GO
911937|T121|Ara-C (Cytarabine), Daunorubicin, Etoposidem, Gemtuzumab Ozogamicin
35803672|T121|Cisplatin and Fluorouracil (CF) and RT
35803672|T121|CF and RT
35803672|T121|Cisplatin, Fluorouracil, Radiation Therapy
35803672|T121|Cisplatin, Fluorouracil Radiation Therapy
35803672|T121|<b>C</b>isplatin, Fluourouracil, Radiation Therapy
35803672|T121|FP and RT
35803672|T121|Fluorouracil, Platinol (Cisplatin), Radiation Therapy
35803672|T121|<b>C</b>isplatin, Fluorouracil, Radiation Therapy
35803673|T121|Fluorouracil, Mitomycin, RT
35803673|T121|Fluorouracil, Mitomycin, Radiation Therapy
35803674|T121|Radiation therapy
35803674|T121|Radiation Therapy
35803674|T121|Involved Field Radiation Therapy
35803675|T121|Non-curative first-line therapy
35803676|T121|Cisplatin and Fluorouracil (CF)
35803676|T121|CF
35803676|T121|FP
35803676|T121|Fluorouracil and Platinol (Cisplatin)
35803676|T121|Cisplatin, Fluorouracil
35803676|T121|Fluorouracil, Platinol (Cisplatin)
35803676|T121|Fluorouracil, Platinol
35803676|T121|Platinol (Cisplatin) and Fluorouracil
35803676|T121|Fluorouracil and Platinol
35802849|T121|mDCF
35802849|T121|modified Docetaxel, Cisplatin, Fluorouracil
35803677|T121|Nivolumab monotherapy
35803678|T121|Pembrolizumab monotherapy
35803678|T121|"<table class=""wikitable"" style=""color:white; background-color:#9e4244"">"
35803678|T121|"<table class=""wikitable"" style=""color:white; background-color:#404040"">"
35803679|T121|Carmustine monotherapy
35803680|T121|CNS cancer surgery
35803681|T121|Lomustine, Vincristine, Prednisone
911920|T121|capmatinib
911920|T121|INC280
911920|T121|Capmatinib
911938|T121|Capmatinib monotherapy
35803682|T121|PCV
35803682|T121|Procarbazine, CCNU, Vincristine
35803682|T121|Procarbazine, CCNU (Lomustine), Vincristine
35803683|T121|RT, then Carmustine
35803684|T121|RT, then Temozolomide
911939|T121|ACP
35803685|T121|Temozolomide, then Temozolomide and RT, then Temozolomide
35803686|T121|Temozolomide and RT
35803686|T121|Temozolomide and Radiation Therapy
35803687|T121|Temozolomide and RT, then Temozolomide
35803688|T121|Bevacizumab monotherapy
35803688|T121|"<table class=""wikitable"" style=""color:white; background-color:#9e4244"">"
35803689|T121|Carboplatin and Bevacizumab
35803690|T121|Cyclophosphamide monotherapy
35803691|T121|Etoposide monotherapy
35803692|T121|Irinotecan monotherapy
911940|T121|PVI
35102014|T121|R-CHOP (Prednisolone)
35102014|T121|Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisolone
35803693|T121|Irinotecan and Bevacizumab
35102013|T121|R-CHOP (Rituximab and hyaluronidase)
35102013|T121|Rituximab and hyaluronidase, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisolone
35803694|T121|Emesis prevention
35102012|T121|R-CHOP-14 (Prednisolone)
35102012|T121|Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisolone every 14 days
35102011|T121|R-MCP (CCNU)
35102011|T121|Rituximab, Methotrexate, CCNU (Lomustine), Procarbazine
35803695|T121|APO
35803695|T121|Adriamycin (Doxorubicin), Prednisone, Oncovin (Vincristine)
35803695|T121|Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone
35803696|T121|BV-CHP
35803696|T121|Brentuximab Vedotin, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Prednisone
35803696|T121|A+CHP
35803696|T121|Adcetris (Brentuximab vedotin), Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Prednisone
35803697|T121|CHOEP-14
35803697|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Etoposide, Prednisone every 14 days
35803697|T121|CHOPE
35803697|T121|VACOP
35803697|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne, Etoposide
35803697|T121|Vepesid (Etoposide), Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Prednisone
35803698|T121|CHOEP-21
35803698|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Etoposide, Prednisone every 21 days
35803698|T121|CHOPE
35803698|T121|VACOP
35803698|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne, Etoposide
35803698|T121|Vepesid (Etoposide), Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Prednisone
35803699|T121|CHOP
35803699|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone
35803699|T121|CHOP-21
35803699|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone every 21 days
35803699|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
35803700|T121|DA-EPOCH
35803700|T121|Dose Adjusted Etoposide, Prednisone, Oncovin (Vincristine), Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin)
35803701|T121|Trimethoprim/Sulfamethoxazole (Bactrim DS)
35803702|T121|Brentuximab vedotin monotherapy
35803703|T121|DHAP
35803703|T121|Dexamethasone, High-dose Ara-C (cytarabine), Platinol (cisplatin)
35803703|T121|Dexamethasone, High-dose Ara-C (Cytarabine), Platinol (Cisplatin)
35803704|T121|GDP
35803704|T121|Gemcitabine, Dexamethasone, Platinol (Cisplatin)
35803705|T121|FluBuCy, then allo HSCT
35803705|T121|FluBuCy
35803706|T121|Altraz
35803707|T121|Anabrez
35803708|T121|Anastraze
35803709|T121|Anastrazol Rontag
35803710|T121|Anastrol
35803711|T121|Arimidex
35803712|T121|Asiolex
35803713|T121|Karomex
35803714|T121|Leprofen
35803715|T121|RUI SI YI
35803716|T121|RUI Ting
35803717|T121|Trozolet
35803718|T121|Trozolite
35803719|T121|FEIBA NF
35803720|T121|Warfarin monotherapy
42542257|T121|enfortumab vedotin-ejfv
42542257|T121|ASG-22CE
42542257|T121|Enfortumab vedotin
42542258|T121|Enfortumab vedotin monotherapy
42542258|T121|"<table class=""wikitable"" style=""color:white; background-color:#9e4244"">"
35803721|T121|Rivaroxaban monotherapy
35803722|T121|ATryn
35803723|T121|Thrombate III
35803724|T121|Atgam
35803725|T121|Lymphoglobuline
35803726|T121|Thymogam
35803727|T121|ATG-Fresenius
35803728|T121|Grafalon
35803729|T121|Thymoglobulin
35803730|T121|Erleada
35803731|T121|Aitan
35803732|T121|Eliquis
35803733|T121|ATG (Horse) and Cyclosporine
35803733|T121|ATG and Cyclosporine
35803733|T121|ATG and CsA
35803733|T121|AntiThymocyte Globulin and Cyclosporine
35803733|T121|AntiThymocyte Globulin and Cyclosporine A
42542259|T121|Enhertu
42542260|T121|DS-8201a
42542260|T121|fam-trastuzumab deruxtecan-nxki
42542260|T121|Trastuzumab deruxtecan
42542261|T121|Fam-trastuzumab deruxtecan monotherapy
35803734|T121|ATG (Horse), Cyclosporine, Eltrombopag
911941|T121|Isa-PD
35803735|T121|ATG (Horse), Cyclosporine, Methylprednisolone
35803736|T121|ATG (Horse), Cyclosporine, G-CSF
35803737|T121|ATG (Horse), Cyclosporine, Sirolimus
35803738|T121|ATG (Rabbit) and Cyclosporine
35803739|T121|Cyclosporine monotherapy
35803741|T121|Eltrombopag monotherapy
35803742|T121|Cinvanti
35803743|T121|Emend
35803744|T121|Emend Trifold
35803745|T121|Acova
35803746|T121|Exembol
35803747|T121|Novastan
35803748|T121|Arsenol
35803749|T121|Arsenox
35803750|T121|Leusenox
35803751|T121|Trisenox
35803752|T121|Asparaginasa
35803753|T121|Chephacardin
35803754|T121|Crasnitin
35803755|T121|Elspar
35803756|T121|Engenase
35803757|T121|Kidrolase
35803758|T121|Laspar
35803759|T121|L Asparaginasa
35803760|T121|L Asparaginasum
35803761|T121|L-Asperone
35803762|T121|L-Ginase
35803763|T121|Leucoginase
35803764|T121|Leunase
35803765|T121|Onconase
35803766|T121|Paronal
35803767|T121|Erwinase
35803768|T121|Erwinaze
35803769|T121|Acard
35803770|T121|Acenterine
35803771|T121|Acesal
35803772|T121|Acesan
35803773|T121|Acetard
35803774|T121|Acetisal
35803775|T121|Acetophen
35803776|T121|Acetosal
35803777|T121|Acetylsalicylsaeure
35803778|T121|Acetylsalicylsyra
35803779|T121|Acetylsalicylsyre
35803780|T121|Acetylsalicylzuur
35803781|T121|Acetylsalisylsyre
35803782|T121|Acetysal
35803783|T121|Acisal
35803784|T121|Actispirine
35803785|T121|Acylpyrin
35803786|T121|Adiprin
35803787|T121|Albyl
35803788|T121|Albyl-Selters
35803789|T121|Albyl Minor
35803790|T121|Anbol
35803791|T121|Ancasal
35803792|T121|Andol
35803793|T121|Angettes
35803794|T121|Anopyrin
35803795|T121|Artria-SR
35803796|T121|Asacard
35803797|T121|Asaferm
35803798|T121|Asaflow
35803799|T121|Asalent
35803800|T121|Asalite
35803801|T121|Asaphen
35803802|T121|Asarid
35803803|T121|Ascardia
35803804|T121|Asdol
35803805|T121|Aspecard
35803740|T121|Aspent
35803806|T121|Aspenter
35803807|T121|Asperan
35803808|T121|Aspergic
35803809|T121|Aspergum
35803810|T121|Aspeter
35803811|T121|Aspilets
35803812|T121|Aspirina-G
35803813|T121|Aspirina
35803814|T121|Aspirine
35803815|T121|Aspirinetas
35803816|T121|Aspirinetta
35803817|T121|Aspirisucre
35803818|T121|Aspirtab
35803819|T121|Aspisol
35803820|T121|Aspocid
35803821|T121|Asprim
35803822|T121|Asprimox ID
35803823|T121|Aspro
35803824|T121|Asrin
35803825|T121|Astrix
35803826|T121|Ataspin
35803827|T121|Avasyl
35803828|T121|Babyprin
35803829|T121|Babypyrin
35803830|T121|Baludon
35803831|T121|Bamycor
35803832|T121|Bamyl
35803833|T121|Bamyl S
35803834|T121|Bayaspirin
35803835|T121|Bayaspirina
35803836|T121|Bestpirin
35803837|T121|Bioplak
35803838|T121|Bokey EMC
35803839|T121|Breoprin
35803840|T121|Bufacyl
35803841|T121|Buferin
35803842|T121|Bufferin
35803843|T121|Cafenol
35803844|T121|Cafiaspirina
35803845|T121|Caprin
35803846|T121|Capsasal
35803847|T121|Cardegic
35803848|T121|Cardioaspirina
35803849|T121|Cardioaspirine
35803850|T121|Cardiopirin
35803851|T121|Cardirene
35803852|T121|Casprium
35803853|T121|Catalgine
35803854|T121|Catalgix
35803855|T121|CC COR
35803856|T121|Cebaspirine
35803857|T121|Cemirit
35803858|T121|Claradin
35803859|T121|Claragine
35803860|T121|Clariprin
35803861|T121|Colfarit
35803862|T121|Colsprin
35803863|T121|Contra-Schmerz ASS
35803864|T121|COR-30
35803865|T121|Coraspin
35803866|T121|Coraspirina
35803867|T121|Corplus
35803868|T121|Corsalbene
35803869|T121|Coryphen
35803870|T121|Delgesic
35803871|T121|Demoprin Novum
35803872|T121|Disperin
35803873|T121|Dispril
35803874|T121|Disprin
35803875|T121|Disprina
35803876|T121|Doloderm
35803877|T121|Doloprin
35803878|T121|Dolorosan
35803879|T121|Draspir
35803880|T121|Dulcipirina
35803881|T121|Dusil
35803882|T121|Easprin
35803883|T121|Ecopirin
35803884|T121|Ecoprin
35803885|T121|Ecosprin
35803886|T121|Ecotrin
35803887|T121|Ecotrin 650
35803888|T121|Ecotrin Maximum Strenght
35803889|T121|Egicalm
35803890|T121|Empirin
35803891|T121|Encaprin
35803892|T121|Encoprin
35803893|T121|Enterosarine
35803894|T121|Entrophen
35803895|T121|Equate Daily
35803896|T121|Fitoaspirin
35803897|T121|Flectadol
35803898|T121|Garaspirine
35803899|T121|Geniol AP
35803900|T121|Geniolito
35803901|T121|Geniol SC
35803902|T121|Geniol SC SIN Cafeina
35803903|T121|Genprin
35803904|T121|Globentyl
35803905|T121|Godamed TAH
35803906|T121|Halfprin
35803907|T121|Herzass
35803908|T121|Hjerdyl
35803909|T121|Hjertealbyl
35803910|T121|Huma ASA
35803911|T121|Hybin
35803912|T121|Junior Asprin
35803913|T121|Jusprin
35803914|T121|Karmyl
35803915|T121|Kilios
35803916|T121|Lasdol
35803917|T121|Levius
35803918|T121|Licyl
35803919|T121|Lisaspin
35803920|T121|LO-Aspirin
35803921|T121|Lowasa
35803922|T121|Lysoprin
35803923|T121|Magnecyl
35803924|T121|Measurin
35803925|T121|Medi-RUB
35803926|T121|Medisyl
35803927|T121|Mejoral Infantil
35803928|T121|Melhoral Infantil
35803929|T121|Metaspirine
35803930|T121|Micristin
35803931|T121|Micropirin
35803932|T121|Migraspirina
35803933|T121|Miniasal
35803934|T121|Minimax
35803935|T121|Naspro
35803936|T121|Nichiaspirin
35803937|T121|Nova-Phase
35803938|T121|Novasen
35803939|T121|Novid
35803940|T121|Pharmacin
35803941|T121|Pharmaspirin
35803942|T121|Phenaspirine
35803943|T121|Platet
35803944|T121|Polopiryna
35803945|T121|Polopiryna S
35803946|T121|Premaspin
35803947|T121|Primaspan
35803948|T121|Quinton
35803949|T121|Remin S
35803950|T121|Reumyl
35803951|T121|Rhodine
35803952|T121|Rhonal
35803953|T121|Rhusal
35803954|T121|Rivasa
35803955|T121|Ronal
35803956|T121|S.R.A.
35803957|T121|SAL-Adult
35803958|T121|Salitison
35803959|T121|Salospir
35803960|T121|Salospir-A
35803961|T121|Saspryl
35803962|T121|Sinaspir
35803963|T121|Solprin
35803964|T121|Solpyron
35803965|T121|Soluble AAC
35803966|T121|Solusprin
35803967|T121|Spren
35803968|T121|Stanback
35803969|T121|Stanback Analgesic
35803970|T121|Supasa
35803971|T121|Tampyrine
35803972|T121|Thomapyrin Akut
35803973|T121|Thrombace NEO
35803974|T121|Thrombo
35803975|T121|Thrombo AS
35803976|T121|Thrombo ASS
35803977|T121|Togal ASS
35803978|T121|Toldex
35803979|T121|Tooprin
35803980|T121|Tromalyt
35803981|T121|Trombyl
35803982|T121|Uniaspirin
35803983|T121|Upsalgina
35803984|T121|Upsarin
35803985|T121|Venopirin
35803986|T121|Winsprin
35803987|T121|Zenaspirin
35803988|T121|Zoprin
35803989|T121|Zorprin
35803990|T121|Aggrenox
35803991|T121|Tecentriq
35803992|T121|Mepron
35803993|T121|Atropen
35803994|T121|Eculizumab monotherapy
42542262|T121|Hemolytic process
911942|T121|Kevadon
35803995|T121|Sirolimus monotherapy
35803996|T121|BCNU/TT
35803996|T121|BCNU (Carmustine), ThioTepa
35803997|T121|BEAC
35803997|T121|BiCNU (Carmustine), Etoposide, Ara-C (Cytarabine), Cyclophosphamide
35803997|T121|Rituximab, BiCNU (Carmustine), Etoposide, Ara-C (Cytarabine), Cyclophosphamide
35803998|T121|BeEAM
35803998|T121|Bendamustine, Etoposide, Ara-C (Cytarabine), Melphalan
35803999|T121|Bortezomib and Melphalan
35803999|T121|Bor-HDM
35803999|T121|Bortezomib, High Dose Melphalan
35804000|T121|Busulfan and Melphalan
35804000|T121|BuMel
911943|T121|Maygace
911944|T121|Megestat
35804001|T121|Bu/TT
35804001|T121|Busulfan, ThioTepa
911945|T121|Anti-BCMA antibody
911946|T121|Megestil
35804002|T121|Bu/TT/Cy
35804002|T121|TBC
35804002|T121|Busulfan, ThioTepa, Cyclophosphamide
35804002|T121|Thiotepa, Busulfan, , Cyclophosphamide
35804002|T121|Thiotepa, Busulfan, Cyclophosphamide
35804003|T121|CBV
35804003|T121|Cyclophosphamide, BiCNU (Carmustine), VP-16 (Etoposide)
35804004|T121|CBV-Mx
35804004|T121|Cyclophosphamide, BiCNU (Carmustine), VP-16 (Etoposide), Mitoxantrone
35804005|T121|CHUT
35804006|T121|CTCb
35804006|T121|Cyclophosphamide, Thiotepa, Carboplatin
911947|T121|Neurosedyn
911948|T121|Niagestin
35804007|T121|Cyclophosphamide, Etoposide, TBI
35804008|T121|FEAM
35804008|T121|Fotemustine, Etoposide, Ara-C (Cytarabine), Melphalan
35804009|T121|LEED
35804009|T121|L-PAM (Melphalan), Endoxan (Cyclophosphamide), Etoposide, Dexamethasone
35804010|T121|Melphalan and TBI
35804010|T121|Melphalan and Total Body Irradiation
35804011|T121|Melphalan monotherapy
35804011|T121|P
35804011|T121|Phenylalanine mustard (Melphalan)
35804011|T121|HDM
35804011|T121|High-Dose Melphalan
911949|T121|Orimentin
35804012|T121|R-BEAM
35804012|T121|Rituximab, BiCNU (Carmustine), Etoposide, Ara-C (Cytarabine), Melphalan
911950|T121|Ovaban
35804013|T121|R-TBI/Cy
35804013|T121|Rituximab, Total, Body, Irradiation, Cyclophosphamide
35804014|T121|TAM6
35804014|T121|Total-body irradiation, Ara-C (Cytarabine), Melphalan
911951|T121|Pallace
35804015|T121|TBI
35804015|T121|Total Body Irradiation
911952|T121|Pantosediv
35804016|T121|Z-BEAM
35804016|T121|Zevalin (Ibritumomab tiuxetan), BiCNU (Carmustine), Etoposide, Ara-C (Cytarabine), Melphalan
35804017|T121|Bendamustine monotherapy
35804018|T121|Doptelet
35804019|T121|Bavencio
35804020|T121|Yescarta
35804021|T121|Inlyta
35804022|T121|Azacitidina
35804023|T121|Azacytin
35804024|T121|Azadine
35804025|T121|Azafect
35804026|T121|Azaplast
35804027|T121|Citaza
35804028|T121|MyAza
35804029|T121|Myelotex
35804030|T121|Vidaza
35804031|T121|Xpreza
35804032|T121|Cyclophosphamide, Daunorubicin, L-Asparaginase, Vincristine, Prednisone
35804033|T121|DOLP
35804033|T121|DVPA
35804033|T121|Daunorubicin, Oncovin (Vincristine), L-Asparaginase, Prednisone
35804033|T121|Daunorubicin, Vincristine, Prednisone, Asparaginase
35804034|T121|Imatinib and Prednisone
35804035|T121|Vincristine and Prednisone
35804035|T121|VP
35804036|T121|Cyclophosphamide, Cytarabine, Mercaptopurine
35804037|T121|Daunorubicin, L-Asparaginase, Vincristine, Prednisone, Imatinib
35804038|T121|L-Asparaginase and Methotrexate
35102010|T121|TH-FEC and H (Docetaxel, SC Trastuzumab)
35102010|T121|TH-FEC and H
35102010|T121|Taxotere (Docetaxel) and Herceptin Hylecta (Trastuzumab and hyaluronidase), followed by Fluorouracil, Epirubicin, Cyclophosphamide, Herceptin Hylecta (Trastuzumab and hyaluronidase)
35102009|T121|FULV (L-Leucovorin)
35102009|T121|5-FU and LevoLeucoVorin
35102008|T121|FOLFIRI (L-Leucovorin)
35102008|T121|L-FOLinic acid, Fluorouracil, IRInotecan
35804040|T121|Cyclophosphamide, Daunorubicin, Vincristine, Prednisone
911953|T121|GSK2857916
911953|T121|belantamab mafodotin-blmf
911953|T121|Belantamab mafodotin
35804041|T121|Pediatric-like GRAALL consolidation
35102007|T121|FOLFIRI and Bevacizumab (L-Leucovorin)
35102007|T121|L-FOLinic acid, Fluorouracil, IRInotecan, Bevacizumab
35102006|T121|FOLFIRI and Cetuximab (L-Leucovorin)
35102006|T121|L-FOLinic acid, Fluorouracil, IRInotecan, Cetuximab
911954|T121|Cisplatin and Bevacizumab
911955|T121|Rodazol
911956|T121|Belantamab mafodotin monotherapy
35804043|T121|Cyclophosphamide, Daunorubicin, L-Asparaginase, Vincristine, Prednisone, Rituximab
35804044|T121|Cytarabine, Idarubicin, Rituximab
35804045|T121|Cyclophosphamide, Idarubicin, Vincristine, Prednisone
35804046|T121|Linker regimen (consolidation)
35102005|T121|FOLFOX 7/sLV5FU2 (L-Leucovorin)
35102005|T121|L-FOLinic acid, Fluorouracil, OXaliplatin alternating with simplified L-LeucoVorin, 5-FU, 2-weekly (every 2 weeks)
35102004|T121|FOLFOX4 (L-Leucovorin)
35102004|T121|L-FOLinic acid, Fluorouracil, OXaliplatin
911957|T121|Sarclisa
911958|T121|Sedalis
911959|T121|Sedoval K17
911960|T121|Single-agent cytotoxic chemotherapy regimen
911961|T121|Single-agent endocrine therapy regimen
911962|T121|Single-agent hypomethylating agent regimen
911963|T121|Single-agent immunotherapy regimen
35804047|T121|Daunorubicin, Pegaspargase, Vincristine, Dexamethasone
35804048|T121|Daunorubicin, Pegaspargase, Vincristine, Prednisone
911964|T121|Single-agent targted therapy regimen
35804049|T121|Hyper-CVAD/MA
35804049|T121|Hyperfractionated Cyclophosphamide, Vincristine, Adriamycin (Doxorubicin), Dexamethasone alternating with Methotrexate, Ara-C (Cytarabine)
911965|T121|Softenon
35804050|T121|Mini-Hyper-CVD/MA and Inotuzumab ozogamicin
35804050|T121|Mini (lower intensity) Hyperfractionated Cyclophosphamide, Vincristine, Dexamethasone alternating with Methotrexate and Ara-C (Cytarabine) and Inotuzumab ozogamicin
911966|T121|Supprelin
35804051|T121|R-Hyper-CVAD/R-MA
35804051|T121|Rituximab, Hyperfractionated Cyclophosphamide, Vincristine, Adriamycin (Doxorubicin), Dexamethasone alternating with Rituximab, Methotrexate, Ara-C (Cytarabine)
35804051|T121|Rituximab, Hyperfractionated Cyclophosphamide, Vincristine, Adriamycin (Doxorubicin), Dexamethasone altenating with Rituximab, Methotrexate, Ara-C (Cytarabine)
911967|T121|FULV and Trimetrexate
35804052|T121|CALGB 8811 regimen
35804053|T121|Mercaptopurine, Methotrexate, WB-XRT
35804054|T121|International ALL Trial
911968|T121|Synovir
35804055|T121|Augmented BFM consolidation
911969|T121|Talimol
35804056|T121|Blinatumomab monotherapy
35804057|T121|Etoposide and TBI, then allo HSCT
35804058|T121|Mercaptopurine, Methotrexate, Vincristine
35804058|T121|BFM HDMTX
35804058|T121|Berlin Frankfurt Muenster High-Dose MTX (Methotrexate) regimen
911970|T121|Tarvacin
911971|T121|Thalido
35804059|T121|Methotrexate and Vincristine
911972|T121|Thalimide
35804060|T121|Augmented Hyper-CVAD and Asparaginase
911973|T121|Thalitero
911974|T121|Thaloma
911975|T121|Blenrep
911976|T121|irbinitinib
911976|T121|ARRY-380
911976|T121|ONT-380
911976|T121|Tucatinib
35804061|T121|CCE
35804061|T121|Clofarabine, Cyclophosphamide, Etoposide
35804062|T121|Daunorubicin, L-Asparaginase, Vincristine, Prednisone
35804063|T121|Hyper-CVAD/MA and Everolimus
35804063|T121|Hyperfractionated Cyclophosphamide, Vincristine, Adriamycin (Doxorubicin), Dexamethasone alternating with Methotrexate, Ara-C (Cytarabine), with Everolimus
35804064|T121|Inotuzumab ozogamicin monotherapy
35804065|T121|Mitoxantrone, Pegaspargase, Vincristine, Dexamethasone
35804066|T121|Tisagenlecleucel monotherapy
911977|T121|Yonsa
35804067|T121|Vincristine liposomal monotherapy
35804068|T121|Non-curative subsequent-line maintenance therapy
35804069|T121|Dasatinib and Prednisone
42542263|T121|Ph-positive B-cell acute lymphoblastic leukemia
35804070|T121|Daunorubicin, Vincristine, Prednisolone, Nilotinib
35804071|T121|Nilotinib-based consolidation
35804072|T121|Hyper-CVAD/MA and Dasatinib
35804072|T121|Hyperfractionated Cyclophosphamide, Vincristine, Adriamycin (Doxorubicin), Dexamethasone alternating with Methorexate and Ara-C (Cytarabine) and Dasatinib
35804073|T121|Hyper-CVAD/MA and Imatinib
35804073|T121|Hyperfractionated Cyclophosphamide, Vincristine, Adriamycin (Doxorubicin), Dexamethasone alternating with Methorexate and Ara-C (Cytarabine) and Imatinib
35102003|T121|Aacidexam
35804074|T121|Hyper-CVAD/MA and Ponatinib
35804074|T121|Hyperfractionated Cyclophosphamide, Vincristine, Adriamycin (Doxorubicin), Dexamethasone alternating with Methorexate and Ara-C (Cytarabine) and Ponatinib
35102002|T121|AALL0232 consolidation
35804075|T121|HAM and Imatinib
35804075|T121|High-dose Ara-C (Cytarabine) and Mitoxantrone and Imatinib
35804076|T121|Imatinib, Vincristine, Dexamethasone
35804077|T121|Cytarabine, Idarubicin, Imatinib
35804078|T121|Imatinib-based consolidation
35804079|T121|Nilotinib monotherapy
35804080|T121|Dasatinib monotherapy
35804081|T121|Dasatinib, Vincristine, Prednisone
35804082|T121|Bosutinib monotherapy
35102001|T121|Abacin
35804083|T121|Imatinib monotherapy
35102000|T121|Abactrim
35804084|T121|Ponatinib monotherapy
35804085|T121|Aminopterin monotherapy
35804086|T121|COMP
35804086|T121|Cyclophosphamide, Oncovin (Vincristine), Methotrexate, Prednisone
911978|T121|daratumumab and hyaluronidase-fihj
911978|T121|Daratumumab and hyaluronidase
35804087|T121|Cyclophosphamide, Doxorubicin, L-Asparaginase, Vincristine, Prednisolone
35804088|T121|Cytarabine, Daunorubicin, L-Asparaginase, Vincristine, Dexamethasone
35804089|T121|Cytarabine, Daunorubicin, L-Asparaginase, Teniposide, Vincristine, Prednisone
911979|T121|Daratumumab and hyaluronidase monotherapy
35101999|T121|Abatrim
911980|T121|Darzalex Faspro
35804090|T121|Doxorubicin, Methotrexate, Vincristine, Prednisone
911981|T121|Daunorubicin, Pegaspargase, Vincristine, Prednisone, Dasatinib
35804091|T121|L-Asparaginase, Vincristine, Dexamethasone
911982|T121|Daunorubicin, Pegaspargase, Vincristine, Prednisone, Imatinib
35804092|T121|L-Asparaginase, Vincristine, Prednisolone
35804092|T121|LVP
35804092|T121|L-asparaginase, Vincristine, Prednisolone
35804093|T121|L-Asparaginase, Vincristine, Prednisone
911983|T121|BTH (Taxotere)
35804094|T121|Mercaptopurine and Prednisone
35804095|T121|Methotrexate monotherapy
35804096|T121|Bacillus Calmette-Guerin (BCG) monotherapy
35804096|T121|"<table class=""wikitable"" style=""color:white; background-color:#9e4244"">"
35804097|T121|Daunorubicin and Prednisone
35804098|T121|Pentostatin monotherapy
35804099|T121|TBI, then auto HSCT
35804100|T121|Dabrafenib and Trametinib
42542264|T121|BRAF-mutated malignancy
35804101|T121|Vemurafenib monotherapy
35804102|T121|TheraCys
35804103|T121|TICE BCG
35804104|T121|Beleodaq
35804105|T121|Camptobell
35804106|T121|Bendamax
35804107|T121|Bendawel
35804108|T121|Bendeka
35804109|T121|Bendit
35804110|T121|Innomustine
35804111|T121|Leuben
35804112|T121|Levact
35804113|T121|Maxtorin
35804114|T121|MyMust
35804115|T121|Purplz
35804116|T121|Ribomustin
35804117|T121|Treakisym
35804039|T121|Treanda
35804118|T121|Xyotin
35804119|T121|Bevyxxa
35804120|T121|Mvasi
35804042|T121|Altuzan
35804121|T121|Avastin
35804122|T121|BevaciRel
35804123|T121|Bevarest
35804124|T121|Bexgratin
35804125|T121|Targretin
35804126|T121|Casodex
35804127|T121|Cosudex
35804128|T121|Calutide
35804129|T121|Kalumid
35804130|T121|Mektovi
35804131|T121|Angiomax
35804132|T121|Angiox
35804133|T121|Local therapy
35804134|T121|Doxorubicin monotherapy
35804134|T121|A
35804134|T121|Adriamycin (Doxorubicin)
35804135|T121|Gemcitabine monotherapy
35804135|T121|"<table class=""wikitable"" style=""color:white; background-color:#9e4244"">"
35804136|T121|Mitomycin monotherapy
35804137|T121|Nephroureterectomy
35804139|T121|Pirarubicin monotherapy
35804140|T121|Thiotepa monotherapy
35804141|T121|Neoadjuvant therapy
35804142|T121|Bladder cancer surgery
35804143|T121|MCV
35804143|T121|CMV
35804143|T121|Methotrexate, Cisplatin, Vinblastine
35804143|T121|Cisplatin, Methotrexate, Vinblastine
35804144|T121|Cisplatin and RT
35804144|T121|Cisplatin and Radiation Therapy
35804145|T121|Cystectomy
35101998|T121|Abditri
35804146|T121|MVAC
35804146|T121|Methotrexate, Vinblastine, Adriamycin (Doxorubicin), Cisplatin
35804146|T121|Methotrexate, Vinblastine, Adriamycin, Cisplatin
35804147|T121|Radical cystectomy
35804148|T121|MVAC, dose-dense
35804148|T121|ddMVAC
35804148|T121|AMVAC
35804148|T121|dose-dense Methotrexate, Vinblastine, Adriamycin (Doxorubicin), Cisplatin
35804148|T121|Accelerated Methotrexate, Vinblastine, Adriamycin (Doxorubicin), Cisplatin
35804148|T121|dose-dense Methotrexate, Vinblastine, Adriamycin, Cisplatin
35804149|T121|Radical cystectomy with bilateral lymphadenectomy
35804150|T121|No neoadjuvant therapy
35804151|T121|Cisplatin, Paclitaxel, RT
35804151|T121|Cisplatin, Paclitaxel, Radiation Therapy
35804151|T121|TP and RT
35804151|T121|Taxol (Paclitaxel), Platinol (Cisplatin), Radiation Therapy
35804151|T121|CP and RT
35804152|T121|Gemcitabine and RT
35804152|T121|Gemcitabine and Radiation Therapy
35804153|T121|Paclitaxel and RT
35804153|T121|Paclitaxel and Radiation Therapy
35804154|T121|PGC
35804154|T121|PCG
35804154|T121|Paclitaxel, Gemcitabine, Cisplatin
35804154|T121|Paclitaxel, Cisplatin, Gemcitabine
35804155|T121|Cisplatin and Methotrexate
35101997|T121|Abetrim
911984|T121|Camrelizumab monotherapy
35804138|T121|Atezolizumab monotherapy
35804156|T121|Carboplatin and Gemcitabine (GCb)
35804156|T121|GCb
35804156|T121|Gemcitabine and Carboplatin
35804156|T121|GC
35804156|T121|GCa
35804156|T121|CG
35804156|T121|Carboplatin and Gemcitabine
35804157|T121|CISCA
35804157|T121|CISplatin, Cyclophosphamide, Adriamycin (Doxorubicin)
911985|T121|Docetaxel and Pertuzumab
35804158|T121|Gemcitabine and Paclitaxel
35804158|T121|GP
35804158|T121|GT
35804158|T121|PG
35804158|T121|Gemcitabine and Taxol (Paclitaxel)
35804158|T121|Paclitaxel and Gemcitabine
35804159|T121|Avelumab monotherapy
35804160|T121|Antihistamines
35804162|T121|Docetaxel monotherapy
35804162|T121|T
35804162|T121|Taxotere (Docetaxel)
35804162|T121|dT
35804162|T121|"<div class=""toccolours"" style=""background-color:#eeeeee"">"
35804162|T121|doceTaxel
35804162|T121|"<table class=""wikitable"" style=""color:white; background-color:#9e4244"">"
911986|T121|Encorafenib monotherapy
35804163|T121|Docetaxel and Ramucirumab
35804164|T121|Durvalumab monotherapy
35804165|T121|Erdafitinib monotherapy
911987|T121|Carboplatin, Pegylated liposomal doxorubicin, Bevacizumab
35804166|T121|Paclitaxel monotherapy
35804166|T121|"<table class=""wikitable"" style=""color:white; background-color:#9e4244"">"
35804166|T121|T
35804166|T121|wP
35804166|T121|Taxol (Paclitaxel)
35804166|T121|weekly Paclitaxel
35804167|T121|Paclitaxel, nanoparticle albumin-bound monotherapy
35804168|T121|Pemetrexed monotherapy
35804169|T121|Vinflunine monotherapy
35804170|T121|Tagraxofusp monotherapy
35804171|T121|Blenoxane
35804172|T121|Bleo
35804173|T121|Bleocin
35804174|T121|Bleocip
35804175|T121|Bleopar
35804176|T121|Bleowel
35804177|T121|Blincyto
35804178|T121|Denosumab monotherapy
35804179|T121|Biocure
35804180|T121|Borater
35804181|T121|Bortecad
35804182|T121|Bortemib
35804183|T121|Bortenat
35804184|T121|Bortetrust
35804185|T121|Bortrac
35804186|T121|Borvex
35804187|T121|Borviz
35804188|T121|Botepar
35804189|T121|Bromadene
35804190|T121|Egybort
35804191|T121|Mibor
35804192|T121|Myezom
35804193|T121|Norvelzo
35804194|T121|Ortez
35804195|T121|Velcade
35804161|T121|Zomib
35804196|T121|Zuricade
35804197|T121|Bosulif
35804198|T121|Brachytherapy
35804199|T121|Cyclophosphamide and Doxorubicin (AC)
35804199|T121|AC
35804199|T121|Adriamycin (Doxorubicin) and Cyclophosphamide
35804199|T121|CA
35804199|T121|Cyclophosphamide and Adriamycin (Doxorubicin)
35804200|T121|Neratinib and Paclitaxel
35804201|T121|Paclitaxel and Trastuzumab (TH)
35804201|T121|TH
35804201|T121|T-T
35804201|T121|Taxol (Paclitaxel) and Herceptin (Trastuzumab)
35804201|T121|Taxol (Paclitaxel) and Trastuzumab
35804201|T121| PH
35804201|T121|Paclitaxel and Herceptin (Trastuzumab)
35804201|T121|Taxol (Paclitaxel), Herceptin (Trastuzumab)
35804201|T121|Trastuzumab, Paclitaxel
35804202|T121|Breast cancer surgery
35804203|T121|THL (Paclitaxel)
35804203|T121|THL
35804203|T121|Taxol (Paclitaxel), Herceptin (Trastuzumab), Lapatinib
35804204|T121|Lapatinib and Paclitaxel (TL)
35804204|T121|TL
35804204|T121|Taxol (Paclitaxel) and Lapatinib
35804205|T121|Paclitaxel monotherapy, weekly
35804205|T121|T
35804205|T121|P
35804205|T121|pT
35804205|T121|wP
35804205|T121|wT
35804205|T121|Taxol (Paclitaxel)
35804205|T121|pacliTaxel
35804205|T121|weekly Paclitaxel
35804205|T121|weekly Taxol (Paclitaxel)
911988|T121|FEC and HP
35804206|T121|Cyclophosphamide and Doxorubicin (AC) and Bevacizumab
35804206|T121|AC and Bevacizumab
35804206|T121|Adriamycin (Doxorubicin), Cyclophosphamide, Bevacizumab
35804207|T121|Docetaxel and Bevacizumab
35804208|T121|Dose-dense Cyclophosphamide and Doxorubicin (ddAC)
35804208|T121|ddAC
35804208|T121|dose-dense Adriamycin (Doxorubicin) and Cyclophosphamide
35804209|T121|Paclitaxel monotherapy, dose-dense (q2wk)
35804209|T121|ddT
35804209|T121|dose-dense Taxol (Paclitaxel)
35804209|T121|ddP
35804209|T121|dose-dense Paclitaxel
35101996|T121|Acetato DE Dexametasona
35804210|T121|Docetaxel and Epirubicin (DE)
35804210|T121|DE
35804210|T121|ED
35804210|T121|ET
35804210|T121|Docetaxel and Epirubicin
35804210|T121|Epirubicin and Taxotere (Docetaxel)
35101995|T121|Acetazona
35804211|T121|Cyclophosphamide and Epirubicin (EC)
35804211|T121|EC
35804211|T121|Epirubicin and Cyclophosphamide
35804212|T121|FEC
35804212|T121|CEF
35804212|T121|Fluorouracil, Epirubicin, Cyclophosphamide
35804212|T121|Cyclophosphamide, Epirubicin, Fluorouracil
911989|T121|Cisplatin, Pemetrexed, RT
35804213|T121|DI EC
35804213|T121|Dose-Intense Epirubicin and Cyclophosphamide
35804214|T121|EDC
35804214|T121|Epirubicin, Docetaxel, Capecitabine
35804215|T121|Epirubicin and Paclitaxel (EP)
35804215|T121|ET
35804215|T121|Epirubicin and Taxol (Paclitaxel)
35804216|T121|FAC
35804216|T121|CAF
35804216|T121|Fluorouracil, Adriamycin (Doxorubicin), Cyclophosphamide
35804216|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Fluorouracil
35804216|T121|AFC
35804216|T121|Adriamycin (Doxorubicin), Fluorouracil, Cyclophosphamide
911990|T121|LGD1057
911990|T121|ALRT1057
911990|T121|Alitretinoin
911991|T121|Acetazolamide
35804217|T121|THP (Docetaxel)
35804217|T121|THP
35804217|T121|"<div class=""toccolours"" style=""background-color:#eeeeee"">"
35804217|T121|Taxotere (Docetaxel), Herceptin (Trastuzumab), Pertuzumab
911992|T121|Cobimetinib, Vemurafenib, Atezolizumab
35101994|T121|Acolon
35804218|T121|PET
35804218|T121|Platinol (Cisplatin), Epirubicin, Taxol (Paclitaxel)
35804219|T121|TAC (Docetaxel)
35804219|T121|TAC
35804219|T121|ATC
35804219|T121|Taxotere (Docetaxel), Adriamycin (Doxorubicin), Cyclophosphamide
35804219|T121|Adriamycin (Doxorubicin), Taxotere (Docetaxel), Cyclophosphamide
35804219|T121|Adriamycin (Doxorubicin), Cyclophosphamide, Taxotere (Docetaxel)
35804220|T121|Docetaxel and Trastuzumab (TH)
35804220|T121|TH
35804220|T121|DH
35804220|T121|"<div class=""toccolours"" style=""background-color:#eeeeee"">"
35804220|T121|Taxotere (Docetaxel) and Herceptin (Trastuzumab)
35804220|T121|Docetaxel and Herceptin (Trastuzumab)
35804220|T121|HT
35804220|T121|H+D
35804220|T121|Herceptin (Trastuzumab) and Taxotere (Docetaxel)
35804220|T121|Herceptin (Trastuzumab) and Docetaxel
35804221|T121|Tamoxifen monotherapy
35804222|T121|Trastuzumab monotherapy
35804223|T121|Paclitaxel monotherapy, q3wk
35804223|T121|T
35804223|T121|P
35804223|T121|pT
35804223|T121|Taxol (Paclitaxel)
35804223|T121|pacliTaxel
35804224|T121|CMF
35804224|T121|Cyclophosphamide, Methotrexate, Fluorouracil
35804224|T121|Cyclophosphamide, Methotrexate, 5-Fluorouracil
35804225|T121|THP (Taxol)
35101993|T121|Actrim
35804226|T121|Doxorubicin and Paclitaxel (AT)
35804226|T121|AT
35804226|T121|Adriamycin (Doxorubicin) and Taxol (Paclitaxel)
35804227|T121|Capecitabine monotherapy
35804227|T121|C
35804227|T121|X
35804227|T121|Xeloda (Capecitabine)
35804228|T121|Epirubicin monotherapy
35804228|T121|E
35804229|T121|Mastectomy
911993|T121|Dara-RVd
911993|T121|D-RVd
911993|T121|Daratumumab, Revlimid (Lenalidomide), Velcade (Bortezomib), Dexamethasone
911994|T121|Dara-Kd
911994|T121|D-Kd
911994|T121|KdD
911994|T121|Daratumumab, Kyprolis (Carfilzomib), low-dose dexamethasone
911994|T121|Kyprolis (Carfilzomib), low-dose dexamethasone, Daratumumab
35804231|T121|CMFT
35804231|T121|Cyclophosphamide, Methotrexate, Fluorouracil, Tamoxifen
35804232|T121|Cyclophosphamide and Docetaxel (TC)
35804232|T121|TC
35804232|T121|Taxotere (Docetaxel) and Cyclophosphamide
35804232|T121|Docetaxel and Cyclophosphamide
35804233|T121|Dose-dense Doxorubicin monotherapy
35804233|T121|ddA
35804233|T121|dose-dense Adriamycin (Doxorubicin)
35101992|T121|Aditrim
35804234|T121|ddTH (Taxol)
35804235|T121|Dose-dense Cyclophosphamide monotherapy
35804235|T121|ddC
35804235|T121|dose-dense Cyclophosphamide
35804236|T121|Dose-dense Cyclophosphamide and Epirubicin (ddEC)
35804236|T121|ddEC
35804236|T121|dose-dense Epirubicin and Cyclophosphamide
35804237|T121|Dose-dense FEC
35804230|T121|ddTH (Taxotere)
35804238|T121|Dose-dense Docetaxel monotherapy
35804238|T121|ddT
35804238|T121|ddD
35804238|T121|dose-dense Taxotere (Docetaxel)
35804238|T121|dose-dense Docetaxel
35101991|T121|Adlone
35101929|T121|Adrecort
35101928|T121|Adrekon
35101927|T121|Adrenol
35101926|T121|Adriamycine
35804239|T121|iddEPC
35804239|T121|intense dose-dense Epirubicin, Paclitaxel, Cyclophosphamide
35804239|T121|IDD-ETC
35804239|T121|Intense Dose-Dense Epirubicin, Taxol (Paclitaxel), Cyclophosphamide
35101925|T121|Adronat
35101924|T121|Adtrim
35804240|T121|Goserelin and Tamoxifen
35101923|T121|Advaferon
35101922|T121|Advantan
35804241|T121|Vinorelbine monotherapy
35804241|T121|V
35804242|T121|Vinorelbine and Trastuzumab (VH)
35804242|T121|VH
35804242|T121|Vinorelbine and Herceptin (Trastuzumab)
35804243|T121|Lapatinib and Trastuzumab
35804243|T121|L+T
35101921|T121|Adventan
35101920|T121|Aeroseb-DEX
35101919|T121|Afpred Forte-Dexa
35804244|T121|Docetaxel and Doxorubicin (AT)
35804244|T121|AT
35804244|T121|AD
35804244|T121|Adriamycin (Doxorubicin) and Taxotere (Docetaxel)
35804244|T121|Adriamycin (Doxorubicin) and Docetaxel
911995|T121|Durvalumab and Tremelimumab
35804245|T121|Capecitabine and Bevacizumab
35804245|T121|CB
35804245|T121|CAP-B
35804245|T121|CAPecitabine and Bevacizumab
35804246|T121|Capecitabine and Docetaxel (TX)
35804246|T121|Taxotere (Docetaxel) and Xeloda (Capecitabine)
35804246|T121|CD
35804246|T121|Capecitabine and Docetaxel
35804246|T121|XT
35804246|T121|Xeloda (Capecitabine) and Taxotere (Docetaxel)
35804246|T121|Docetaxel and Capecitabine
35804247|T121|Capecitabine and Paclitaxel
35804247|T121|Taxol (Paclitaxel), Xeloda (Capecitabine)
35804248|T121|Capecitabine and Paclitaxel, nanoparticle albumin-bound
35804249|T121|Pegylated liposomal doxorubicin monotherapy
35804249|T121|Pegylated Liposomal Doxorubicin
35804250|T121|Cyclophosphamide and Epirubicin (EC) and Bevacizumab
35804250|T121|EC and Bevacizumab
35804250|T121|Epirubicin, Cyclophosphamide, Bevacizumab
35804251|T121|Epirubicin and Vinorelbine
911996|T121|Cyclophosphamide and Epirubicin (EC) and Pembrolizumab
911996|T121|EC and Pembrolizumab
911996|T121|Epirubicin, Cyclophosphamide, Pembrolizumab
35804252|T121|FAC and Bevacizumab
35804252|T121|Fluorouracil, Adriamycin (Doxorubicin), Cyclophosphamide, Bevacizumab
911997|T121|Emapalumab and Dexamethasone
911998|T121|Encorafenib and Cetuximab
35804253|T121|FEC and Bevacizumab
35804253|T121|Fluorouracil, Epirubicin, Cyclophosphamide, Bevacizumab
35804254|T121|Cyclophosphamide and Non-pegylated liposomal doxorubicin (MC)
35804254|T121|MC
35804254|T121|Myocet (non-pegylated liposomal doxorubicin) and Cyclophosphamide
35101918|T121|Aidbone
35804255|T121|Paclitaxel and Bevacizumab
35804256|T121|Paclitaxel, nanoparticle albumin-bound and Bevacizumab
35804257|T121|S-1 monotherapy
35804258|T121|Abemaciclib monotherapy
35804259|T121|Capecitabine and Ixabepilone
35804259|T121|XI
35804259|T121|Xeloda (Capecitabine) and Ixabepilone
35804260|T121|Cisplatin and Vinorelbine (CVb)
35804260|T121|CVb
35804260|T121|VC
35804260|T121|Vinorelbine, Cisplatin
35804260|T121|CV
35804260|T121|NP
35804260|T121|PV
35804260|T121|Navelbine (Vinorelbine) and Platinol (Cisplatin)
35804260|T121|Platinol (Cisplatin) and Vinorelbine
35804260|T121|Vinorelbine and Cisplatin
35101917|T121|AK-DEX
911999|T121|AiRuiKa
35804261|T121|Doxorubicin and Bevacizumab
35804262|T121|Non-pegylated liposomal doxorubicin monotherapy
35804262|T121|Non-Pegylated Liposomal Doxorubicin
35804263|T121|Non-pegylated liposomal doxorubicin and Bevacizumab
35804263|T121|NPLD and Bev
35804263|T121|Non-Pegylated Liposomal Doxorubicin and Bevacizumab
35804264|T121|Pegylated liposomal doxorubicin and Bevacizumab
35804264|T121|PLD and Bev
35804264|T121|Pegylated Liposomal Doxorubicin and Bevacizumab
35804265|T121|Eribulin monotherapy
35804266|T121|Gemcitabine and Bevacizumab
35804267|T121|Ixabepilone monotherapy
35804268|T121|Vinorelbine and Bevacizumab
35804269|T121|Olaparib monotherapy
35804269|T121|"<table class=""wikitable"" style=""color:white; background-color:#9e4244"">"
42542265|T121|BRCA-mutated Breast cancer
35804270|T121|Talazoparib monotherapy
35804271|T121|Anastrozole monotherapy
42542266|T121|ER-positive Breast cancer
35804272|T121|Anastrozole and Goserelin
35804273|T121|Letrozole monotherapy
35101916|T121|Aksotran
35804274|T121|Exemestane monotherapy
35804275|T121|Bilateral oophorectomy
35804276|T121|Goserelin monotherapy
912000|T121|Alizapride
35804277|T121|Leuprolide monotherapy
35804278|T121|Tamoxifen and OFS
35804279|T121|Toremifene monotherapy
35804280|T121|Abemaciclib and Anastrozole
35804281|T121|Abemaciclib and Letrozole
35804282|T121|Anastrozole and Fulvestrant
35804283|T121|Anastrozole, Goserelin, Ribociclib
35804284|T121|Fulvestrant monotherapy
35804285|T121|Fulvestrant and Ribociclib
35101915|T121|Albrotran
35101914|T121|Albutrim
35804286|T121|Letrozole and Bevacizumab
35804287|T121|Letrozole and Palbociclib
35804288|T121|Letrozole and Ribociclib
35804289|T121|Goserelin, Ribociclib, Tamoxifen
35101913|T121|Alcorim-F
35101912|T121|Alcot
35101911|T121|Aldocumar
35101910|T121|Aldren
35101909|T121|Aldron
35101908|T121|Aldronac
35101907|T121|Alecast
35101906|T121|Alemax
35101905|T121|Alenat
35804290|T121|Tamoxifen and Prednisolone
35101904|T121|Alenato
35804291|T121|Anastrozole and Trastuzumab
35804292|T121|Lapatinib and Letrozole
35804293|T121|Lapatinib, Letrozole, Trastuzumab
35804294|T121|Abemaciclib and Fulvestrant
35101903|T121|Alenbon
35101902|T121|Alencar
35101901|T121|Alend
42542267|T121|Bilateral adrenalectomy
35101900|T121|Alendene
35101899|T121|Alendex
35101898|T121|Alendil
35804295|T121|Everolimus and Exemestane
35101897|T121|Alendomax
35101896|T121|Alendon
35804296|T121|Everolimus and Tamoxifen
35101895|T121|Alendor
35101894|T121|Alendra 7
35101893|T121|Alendral
35101892|T121|Alendrate
35101891|T121|Alendrin
35101890|T121|Alendro
35101889|T121|Alendromax
35804297|T121|Fulvestrant and Palbociclib
35101888|T121|Alendron
35101887|T121|Alendronat
35101886|T121|Alendronato
35804298|T121|ECH
35804298|T121|Epirubicin, Cyclophosphamide, Herceptin (Trastuzumab)
42542268|T121|HER2-positive Breast cancer
35101885|T121|Alendronhexal
35101884|T121|Alendroninezr
35804299|T121|FEC and H
35804300|T121|TCHP (Docetaxel)
35804300|T121|TCHP
35804300|T121|Taxotere (Docetaxel), Carboplatin, Herceptin (Trastuzumab), Pertuzumab
35101883|T121|Alendroninezuur
35101882|T121|Alendronsaeure
35101881|T121|Alendronstad
35101880|T121|Alendros
35101879|T121|Alenmax
35804301|T121|T-DM1 monotherapy
35804302|T121|T-DM1 and ET
35804302|T121|Trastuzumab-DM1 (Trastuzumab emtansine) and Endocrine Therapy
35804303|T121|GnRH agonists
35804304|T121|Aromatase inhibitors
35804305|T121|Trastuzumab and ET
35804305|T121|Trastuzumab and Endocrine Therapy
35804306|T121|Neratinib monotherapy
35101878|T121|Alenost
35101877|T121|Alent
35804307|T121|TCH (Docetaxel, Carboplatin)
35804307|T121|Taxotere (Docetaxel), Carboplatin, Herceptin (Trastuzumab)
35804308|T121|TCH (Docetaxel, Cyclophosphamide)
35804308|T121|Taxotere, Cyclophosphamide, Herceptin
35101876|T121|Alentop
35101875|T121|Alergolon
35804309|T121|ACH
35804309|T121|Adriamycin (Doxorubicin), Cyclophosphamide, Herceptin (Trastuzumab)
35804310|T121|Capecitabine, Bevacizumab, Trastuzumab
35804311|T121|Capecitabine and Lapatinib
35804312|T121|Capecitabine and Trastuzumab (XH)
35804312|T121|XH
35804312|T121|Xeloda (Capecitabine) and Herceptin
35804313|T121|Pertuzumab and T-DM1
35804313|T121|Pertuzumab and Trastuzumab-DM1 (Trastuzumab emtansine)
35101874|T121|Alfaferone
35101873|T121|Alfalyl
35804314|T121|Pertuzumab and Trastuzumab
35804315|T121|TPC
35804315|T121|Taxol (Paclitaxel), Platinol (Cisplatin), Capecitabine
35804316|T121|Capecitabine and Neratinib
35804317|T121|Capecitabine, Pertuzumab, Trastuzumab
35804317|T121|XHP
35804317|T121|Xeloda (Capecitabine), Herceptin (Trastuzumab), Pertuzumab
42542269|T121|triple negative Breast cancer
35804318|T121|Carboplatin and nab-Paclitaxel
35804318|T121|CnP
35804319|T121|Bevacizumab-containing therapy
35804320|T121|nab-Paclitaxel monotherapy
35804321|T121|nab-Paclitaxel and Atezolizumab
35804322|T121|Enzalutamide monotherapy
35804323|T121|CVAP
35804323|T121|VACP
35804323|T121|Cyclophosphamide, Vincristine, Adriamycin (Doxorubicin), Prednisolone
35804323|T121|Vincristine, Adriamycin (Doxorubicin), Cyclophosphamide, Prednisolone
35101872|T121|Aliot
35804324|T121|ACT
35804324|T121|Adriamycin (Doxorubicin), Cyclophosphamide, Tamoxifen
35804325|T121|CAMFP
35804325|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Methotrexate, Fluorouracil, Prednisone
35804326|T121|Lumpectomy
35804327|T121|CEF/CMF
35804327|T121|Cyclophosphamide, Epirubicin, Fluorouracil alternating with Cyclophosphamide, Methotrexate, Fluorouracil
35804328|T121|CFP
35804328|T121|Cyclophosphamide, Fluorouracil, Prednisone
35804329|T121|CFP and Oophorectomy
35804329|T121|Cyclophosphamide, Fluorouracil, Prednisone and Bilateral Oophorectomy
35804330|T121|CMFL
35804330|T121|Cyclophosphamide, Methotrexate, Fluorouracil, Leucovorin (Folinic acid)
35804331|T121|CMFP
35804331|T121|Cyclophosphamide, Methotrexate, Fluorouracil, Prednisone
35804332|T121|Modified radical mastectomy
35804333|T121|Total mastectomy with low axillary-node dissection
35804334|T121|CMFPT
35804334|T121|Cyclophosphamide, Methotrexate, Fluorouracil, Prednisone, Tamoxifen
35804335|T121|CMFVP
35804335|T121|Cyclophosphamide, Methotrexate, Fluorouracil, Vincristine, Prednisone
35804335|T121|COMFP
35804335|T121|CFPMV
35804335|T121|Cyclophosphamide, Oncovin (Vincristine), Methotrexate, Fluorouracil, Prednisone
35804335|T121|Cyclophosphamide, Fluorouracil, Prednisone, Methotrexate, Vincristine
35804336|T121|CPB
35804336|T121|Cyclophosphamide, Platinol (Cisplatin), BCNU (Carmustine)
35804337|T121|CTCb, then auto HSCT
35804338|T121|ECT
35804338|T121|Epirubicin, Cyclophosphamide, Thiotepa
35804339|T121|FAC and BCG
35804339|T121|Fluorouracil, Adriamycin (Doxorubicin), Cyclophosphamide, BCG
35804340|T121|FNC
35804340|T121|Fluorouracil, Novantrone (Mitoxantrone), Cyclophosphamide
35804340|T121|Cyclophosphamide, Novantrone (Mitoxantrone), Fluorouracil
35804341|T121|Levamisole monotherapy
35804342|T121|MF
35101871|T121|Allenmax
35101870|T121|Allibac
35804343|T121|Methotrexate and Vinblastine (MV)
35804344|T121|Oophorectomy
35804345|T121|PAF
35804345|T121|Phenylalanine mustard (Melphalan), Adriamycin (Doxorubicin), Fluorouracil
35804346|T121|PF
35804346|T121|Phenylalanine mustard (Melphalan) and Fluorouracil
35804347|T121|PFT
35804347|T121|Phenylalanine mustard (Melphalan), 5-Fluorouracil, Tamoxifen
35804348|T121|PT
35804348|T121|Prednisone and Tamoxifen
35804349|T121|TMF
35804349|T121|Thiotepa, Methotrexate, Fluorouracil
35804350|T121|Aminoglutethimide monotherapy
35804351|T121|CAMF
35804351|T121|AFCM
35804351|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Methotrexate, Fluorouracil
35804351|T121|Adriamycin (Doxorubicin), Fluorouracil, Cyclophosphamide, Methotrexate
35804352|T121|CAF and MPA
35804352|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Fluorouracil, MedroxyProgesterone Acetate
35804353|T121|Chlorambucil and Prednisolone
35804354|T121|CHUT, then auto HSCT
35804355|T121|CMFV
35804355|T121|CVMF
35804355|T121|Cyclophosphamide, Methotrexate, Fluorouracil, Vinblastine
35804355|T121|Cyclophosphamide, Vinblastine, Methotrexate, Fluorouracil
35804356|T121|DES monotherapy
35101869|T121|Alont
35804357|T121|Estradiol monotherapy
35804358|T121|Fluoxymesterone monotherapy
35101868|T121|Alovell
35804359|T121|Formestane monotherapy
35101867|T121|BYL719
35101867|T121|Alpelisib
35804360|T121|Medroxyprogesterone monotherapy
42542270|T121|Padcev
35101866|T121|Alpelisib and Fulvestrant
35101865|T121|Alpermell
35101864|T121|Alquimid
35804361|T121|Megestrol monotherapy
35804362|T121|Methotrexate and Thiotepa
35804363|T121|Mitoxantrone monotherapy
35804364|T121|TAD (Tamoxifen)
35804364|T121|Tamoxifen, Aminoglutethimide, Danazol
35804365|T121|VAC (Adriamycin)
35804366|T121|VAP
35804366|T121|Vincristine, Adriamycin (Doxorubicin), Prednisolone
35804367|T121|Adcetris
35804368|T121|Alunbrig
35804369|T121|COP
35804370|T121|COPADM
35804370|T121|Cyclophosphamide, Oncovin (Vincristine), Prednisone, ADriamycin (Doxorubicin), Methotrexate
35804371|T121|R-COPADM
35804371|T121|Rituximab, Cyclophosphamide, Oncovin (Vincristine), Prednisone, ADriamycin (Doxorubicin), Methotrexate
35804372|T121|BASIC
35804372|T121|Brief, Anthracycline-Sparing, Intensive Cyclophosphamide
35804373|T121|CALGB 10-002 regimen
35804374|T121|CODOX-M
35804374|T121|Cyclophosphamide, Oncovin (Vincristine), DOXorubicin, Methotrexate
35804374|T121|Cyclophosphamide, Oncovin, DOXorubicin, Methotrexate
35804375|T121|CODOX-M/IVAC
35804375|T121|Cyclophosphamide, Oncovin (Vincristine), DOXorubicin, Methotrexate alternating with Ifosfamide, Vepesid (Etoposide), Ara-C (Cytarabine)
35804375|T121|Cyclophosphamide, Oncovin, DOXorubicin, Methotrexate alternating with Ifosfamide, Vepesid (etoposide), Ara-C (cytarabine)
35804376|T121|COPAD
35804376|T121|Cyclophosphamide, Oncovin (Vincristine), Prednisone, ADriamycin (Doxorubicin)
35804377|T121|Cytarabine and Methotrexate (CYM)
35804377|T121|CYtarabine, Methotrexate
35804377|T121|CYtarabine and Methotrexate
35804378|T121|DA-R-EPOCH
35804378|T121|Dose Adjusted Rituximab, Etoposide, Prednisone, Oncovin (Vincristine), Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin)
35804379|T121|GMALL-R
35804379|T121|German Multicenter Study Group for the Treatment of Adult Acute Lymphoblastic Leukemia, Rituximab
35804380|T121|R-CODOX-M
35804380|T121|Rituximab, Cyclophosphamide, Oncovin (Vincristine), DOXorubicin, Methotrexate
35804381|T121|R-CODOX-M/R-IVAC
35804381|T121|Rituximab, Cyclophosphamide, Oncovin (Vincristine), DOXorubicin, Methotrexate alternating with Rituximab, Ifosfamide, Vepesid (etoposide), Ara-C (Cytarabine)
35804381|T121|Rituximab, Cyclophosphamide, Oncovin (Vincristine), DOXorubicin, Methotrexate alternating with Rituximab, Ifosfamide, Vepesid (Etoposide), Ara-C (Cytarabine)
35804382|T121|R-CODOX-M (Pegylated liposomal doxorubicin substituted)
35804382|T121|Rituximab, Cyclophosphamide, Oncovin (Vincristine), DOXil (Pegylated liposomal doxorubicin), Methotrexate
35804383|T121|R-CODOX-M/R-IVAC (Pegylated liposomal doxorubicin substituted)
35804383|T121|Rituximab, Cyclophosphamide, Oncovin (Vincristine), DOXil (Pegylated liposomal doxorubicin), Methotrexate alternating with Rituximab, Ifosfamide, Vepesid (Etoposide), Ara-C (Cytarabine)
35804384|T121|Fluoroquinolone
35804385|T121|COPAD/CYVE
35804385|T121|Cyclophosphamide, Oncovin (Vincristine), Prednisone, ADriamycin (Doxorubicin) alternating with CYtarabine, VEpesid (Etoposide)
35804386|T121|Busulfex
35804387|T121|Myleran
35804388|T121|Dexamethasone monotherapy
35804389|T121|Dexamethasone and WBRT
35804390|T121|Alectinib monotherapy
35101863|T121|Altrim
35804391|T121|Ceritinib monotherapy
35804392|T121|Afatinib monotherapy
35804393|T121|Icotinib monotherapy
35804394|T121|Osimertinib monotherapy
912001|T121|Amonafide
35804395|T121|IT Cytarabine and Methotrexate
35804396|T121|IT Cytarabine, Methotrexate, Methylprednisolone
35804397|T121|IT Cytarabine, Methotrexate, Prednisone
35804398|T121|IT Cytarabine and WBRT
35804398|T121|Cytarabine and WBRT
35804398|T121|Cytarabine and Whole Brain Radiation Therapy
35804399|T121|IT Methotrexate monotherapy
35804400|T121|IT Methotrexate and Hydrocortisone
35804401|T121|IT Methotrexate and Methylprednisolone
35804402|T121|IT Methotrexate and WBRT
35804402|T121|IntraThecal Methotrexate and Whole Brain Radiation Therapy
35804403|T121|WBRT
35804403|T121|Whole Brain Radiation Therapy
35804404|T121|Mercaptopurine and WBRT
35804404|T121|Mercaptopurine and Whole Brain Radiation Therapy
35804405|T121|IT Cytarabine, Methotrexate, WBRT
35804405|T121|Cytarabine, Methotrexate, WBRT
35804405|T121|Cytarabine, Methotrexate, Whole Brain Radiation Therapy
35804406|T121|R-CHOEP-14
35804406|T121|Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Etoposide, Prednisone, 14-day cycles
35804407|T121|IT Cytarabine monotherapy
35804408|T121|IT Cytarabine liposomal monotherapy
35804409|T121|Upfront therapy
35804410|T121|Whole brain irradiation
35804410|T121|Whole-Brain Radiation Therapy
35804410|T121|PCI
35804410|T121|Prophylactic Cranial Irradiation
35804411|T121|BCNU/TT, then auto HSCT
35804412|T121|Cytarabine, Methotrexate, Rituximab
35804412|T121|R-HD-MTX/ARA-C
35804412|T121|Rituximab, High-Dose MethoTreXate, ARA-C (Cytarabine)
35804413|T121|MATRix
35804413|T121|Methotrexate, Ara-C (Cytarabine), Thiotepa, Rituximab
35804414|T121|Bu/TT, then auto HSCT
35804415|T121|Lomustine, Methotrexate, Procarbazine
35804415|T121|Methotrexate, CCNU (Lomustine), Procarbazine
35804416|T121|Lomustine, Methotrexate, Procarbazine, Methylprednisolone
35804417|T121|Methotrexate, then Cytarabine
35804418|T121|BEAM, then auto HSCT
35804419|T121|Methotrexate, then Cytarabine and Thiotepa
35804420|T121|Methotrexate and Rituximab
35804421|T121|MPV
35804421|T121|Methotrexate, Procarbazine, Vincristine
35804422|T121|MT-R
35804422|T121|Methotrexate, Temozolomide, Rituximab
35804423|T121|MVBP
35804423|T121|Methotrexate, VP16 (Etoposide), BCNU (Carmustine), MethylPrednisolone
35804424|T121|Nordic Regimen, older patients
35804425|T121|Nordic Regimen, younger patients
35804426|T121|R-MCP
35804426|T121|Rituximab, Mitoxantrone, Chlorambucil, Prednisolone
35804427|T121|R-MP
35804427|T121|Rituximab, Methotrexate, Procarbazine
35804428|T121|Procarbazine monotherapy
35804429|T121|R-MPV
35804429|T121|Rituximab, Methotrexate, Procarbazine, Vincristine
35804430|T121|Bu/TT/Cy, then auto HSCT
35804431|T121|Ifosfamide and Methotrexate
35101862|T121|Amazole
35804432|T121|Temsirolimus monotherapy
35804433|T121|Topotecan monotherapy
35804434|T121|Dabrafenib monotherapy
35804435|T121|Ipilimumab and Nivolumab
35804436|T121|Jevtana
35804437|T121|Cometriq is the brand name for cabozantinib's medullary thyroid cancer indication. Cabometyx is the brand name for cabozantinib's renal cell carcinoma indication
35804438|T121|Asparlas
35804439|T121|Kengreal
35804440|T121|Cabita
35804441|T121|Capebin
35804442|T121|Capegard
35804443|T121|Capnat
35804444|T121|Caposib
35804445|T121|Capsy
35804446|T121|Caxeta
35804447|T121|Citabin
35804448|T121|Flagoda
35804449|T121|Naprocap
35804450|T121|Skemca
35804451|T121|Xeloda
35804452|T121|Xlotabin
35804453|T121|Cablivi
35804454|T121|Biocarb
35804455|T121|Biocarbo
35804456|T121|Bioplatinex
35804457|T121|Biovinate
35804458|T121|Blastocarb
35804459|T121|Bonaplatin
35804460|T121|Boplatex
35804461|T121|Carbo
35804462|T121|Carbokem
35804463|T121|Carbomedac
35804464|T121|Carbomerck
35804465|T121|Carboplat
35804466|T121|Carboplatine
35804467|T121|Carboplatino
35804468|T121|Carboplatinum
35804469|T121|Carbosin
35804470|T121|Carbotanil
35804471|T121|Carbotec
35804472|T121|Carbotinol
35804473|T121|Careptin
35804474|T121|Carplan
35804475|T121|Carplanil
35804476|T121|Carpsol
35804477|T121|Crobextin
35804478|T121|Cycloplatin
35804479|T121|Cycloplatinum
35804480|T121|Emorzim
35804481|T121|Erbakar
35804482|T121|Ercar
35804483|T121|Fauldcarbo
35804484|T121|Ifacap
35804485|T121|Kemocarb
35804486|T121|Megaplatin
35804487|T121|Nealorin
35804488|T121|Neocarb
35804489|T121|Neocarbo
35804490|T121|Oncocarb
35804491|T121|Paraplatin
35804492|T121|Paraplatine
35804493|T121|Pharmaplatin
35804494|T121|Platamine CS
35804495|T121|Platinwas
35804496|T121|Ribocarbo
35804497|T121|Tecnocarb
35804498|T121|Vancel
35804499|T121|CBDCA
35804500|T121|Kyprolis
35804501|T121|Becenun
35804502|T121|BiCNU
35804503|T121|Carmubris
35804504|T121|Leucerom
35804505|T121|Nitrourean
35804506|T121|Nitrumon
35804507|T121|Biodel
35804508|T121|Gliadel wafer
35804509|T121|Cagin
35804510|T121|Cancidas
35804511|T121|Capsain
35804512|T121|Caspogin
35804513|T121|Caspoliv
35804514|T121|Casponova
35804515|T121|Guficap
35804516|T121|Kabifungin
35804517|T121|Letocan
35804518|T121|Profung
35804519|T121|Wofungin
35804520|T121|Bortezomib monotherapy
42542271|T121|Tositumomab and I-131 (Bexxar)
35804521|T121|Siltuximab monotherapy
35804522|T121|TCP
35804522|T121|Thalidomide, Cyclophosphamide, Prednisone
35804523|T121|Tocilizumab monotherapy
35804524|T121|Recentin
35804525|T121|Libtayo
35804526|T121|Zykadia
35804527|T121|Cisplatin and Paclitaxel
35804527|T121|PC
35804527|T121|CP
35804527|T121|Paclitaxel and Cisplatin
35804527|T121|Taxol (Paclitaxel) and Platinol (Cisplatin)
35804527|T121|Platinol (Cisplatin) and Taxol (Paclitaxel)
35804528|T121|Cervical cancer surgery
35804529|T121|Radical hysterectomy
35804530|T121|Carboplatin and RT
35804530|T121|Carboplatin and Radiation Therapy
35804531|T121|Hysterectomy
35101861|T121|Amethapred
35804532|T121|Cisplatin and Fluorouracil (CF) and Hydroxyurea, RT
35804532|T121|Cisplatin, Fluorouracil, Hydroxyurea, RT
35804532|T121|Cisplatin, Fluorouracil, Hydroxyurea, Radiation Therapy
35804533|T121|Cisplatin and Gemcitabine (GC) and RT
35804533|T121|Cisplatin, Gemcitabine, RT
35804533|T121|Cisplatin, Gemcitabine, Radiation Therapy
35804534|T121|Fluorouracil and RT
35804534|T121|5-FluouroUracil and Radiation Therapy
35804534|T121|5-FluoroUracil and Radiation Therapy
35804534|T121|Fluorouracil and Radiation Therapy
35804535|T121|Hydroxyurea and RT
35804535|T121|Hydroxyurea and Radiation Therapy
35101860|T121|Amilene
35804536|T121|Carboplatin and Ifosfamide
35804537|T121|Carboplatin monotherapy
35804538|T121|Cisplatin and Ifosfamide
35804539|T121|Cisplatin and Mitomycin
35804540|T121|Cisplatin, Paclitaxel, Bevacizumab
35804540|T121|CP+Bev
35804540|T121|"<table class=""wikitable"" style=""color:black; background-color:#42f584"">"
35804541|T121|Cisplatin and Topotecan
35804541|T121|TC
35804541|T121|CT
35804541|T121|Topotecan and Cisplatin
35804542|T121|Ifosfamide monotherapy
35101859|T121|Amoxazol
35101858|T121|Amoxicillin
35101857|T121|Amtran
35101856|T121|Amtril
35804543|T121|Paclitaxel and Topotecan
35804543|T121|Topotecan, Paclitaxel
35804544|T121|Paclitaxel, Topotecan, Bevacizumab
35804544|T121|TP+Bev
35804544|T121|Topotecan, Paclitaxel, Bevacizumab
35101855|T121|Amumetazon
35804545|T121|FULV
35804545|T121|5-FU and LeucoVorin (Folinic acid)
35804545|T121|5-FU (Fluorouracil) and Folinic Acid
35804545|T121|LV5FU2
35804545|T121|LeucoVorin (Folinic acid) and 5-FU for 2 days
35804545|T121|LeucoVorin and 5-FU, two days out of the month
35804545|T121|simplified LeucoVorin and 5-FU, two days out of the month
35804545|T121|FF
35804545|T121|Fluorouracil and Folinic acid
35804546|T121|Cetrine
35804547|T121|Cetzine
35804548|T121|Glocet
35804549|T121|Piriteze
35804550|T121|Razene
35804551|T121|Zyrtec
35804552|T121|Cetuxim
35804553|T121|Erbitux
35804554|T121|Epidaza
35804555|T121|Chlor-Trimeton
35804556|T121|Piriton
35804557|T121|Capecitabine and Gemcitabine
35804557|T121|GemCap
35804557|T121|Gemcitabine and Capecitabine
35804557|T121|GEM-CAP
35804557|T121|GEMcitabine and CAPecitabine
35804557|T121|CAP-GEM
35804557|T121|CAPecitabine and GEMcitabine
35804558|T121|Gemcitabine, then Fluorouracil and RT, then Gemcitabine
35804559|T121|GemOx
35804559|T121|Gemcitabine and Oxaliplatin
35804559|T121|GEMOX
35804559|T121|GEMcitabine and OXaliplatin
35804559|T121|mGEMOX
35804559|T121|modified GEMcitabine and OXaliplatin
35804559|T121|Gemcitabine, Oxaliplatin
35101854|T121|Anasmol
35804560|T121|Capecitabine and Mitomycin
35804561|T121|Cisplatin and Gemcitabine (GC) and nab-Paclitaxel
35804562|T121|ECF
35804562|T121|Epirubicin, Cisplatin, Fluorouracil
35804563|T121|FELV
35804563|T121|Fluorouracil , Etoposide and LeucoVorin (Folinic acid)
35804563|T121|Fluorouracil , Etoposide, LeucoVorin (Folinic acid)
35804564|T121|FULV and Gemcitabine
35804564|T121|5-FU, LeucoVorin (Folinic acid), Gemcitabine
35804565|T121|Gemcitabine, Cisplatin, S-1
35804565|T121|GCS
35804566|T121|Gemcitabine and Mitomycin
35804567|T121|Gemcitabine and nab-Paclitaxel
35804567|T121|NG
35804567|T121|Nab-Paclitaxel and Gemcitabine
35804567|T121|AG
35804567|T121|Abraxane (nab-Paclitaxel) and Gemcitabine
35804568|T121|GEMOX-B
35804568|T121|GEMcitabine, OXaliplatin, Bevacizumab
35804569|T121|Regorafenib monotherapy
35804570|T121|Bendamustine and Rituximab (BR)
35804570|T121|BR
35804570|T121|Bendamustine, Rituximab
35804570|T121|R-B
35804570|T121|Bendamustine and Rituximab
35804570|T121|Rituximab and Bendamustine
35804570|T121|RB
35804570|T121|Rituximab, Bendamustine
35804571|T121|Cladribine and Cyclophosphamide (CC)
35804571|T121|CC
35804571|T121|Cladribine, Cyclophosphamide
35804572|T121|Chlorambucil and Obinutuzumab (GClb)
35804572|T121|GClb
35804572|T121|GA101 (Obinutuzumab) and Chlorambucil
912002|T121|Amoxicillin and PPI
35804573|T121|Chlorambucil and Ofatumumab
35804574|T121|Chlorambucil and Rituximab (RClb)
35804574|T121|RClb
35804574|T121|CLB-R
35804574|T121|Rituximab and Chlorambucil
35804574|T121|ChLoramBucil and Rituximab
35804575|T121|CMC
35804575|T121|Cladribine, Mitoxantrone, Cyclophosphamide
35804576|T121|FCA
35804576|T121|FCCam
35804576|T121|Fludarabine, Cyclophosphamide, Alemtuzumab
35804576|T121|Fludarabine, Cyclophosphamide, Campath (Alemtuzumab)
35804577|T121|FCM
35804577|T121|Fludarabine, Cyclophosphamide, Mitoxantrone
35804578|T121|PCP prophylaxis
35804579|T121|Hematopoietic growth factors
912003|T121|Amoxicillin, Clarithromycin, PPI, Bismuth
912004|T121|Ampicillin
35804580|T121|Fludarabine and Alemtuzumab
35804580|T121|Fludarabine and Campath (Alemtuzumab)
35804581|T121|Ibrutinib monotherapy
35804582|T121|Ibrutinib and Obinutuzumab
35804583|T121|Obinutuzumab monotherapy
912005|T121|Ampicillin and PPI
35804584|T121|Alemtuzumab and Methylprednisolone
35804585|T121|Bendamustine and Obinutuzumab
35804585|T121|G-B
35804585|T121|Gazyva (Obinutuzumab), Bendamustine
35804585|T121|Gazyva (Obinutuzumab) and Bendamustine
35804586|T121|Antivirals
35804587|T121|CFAR
35804587|T121|Cyclophosphamide, Fludarabine, Alemtuzumab, Rituximab
35804588|T121|G-FC
35804588|T121|Gazyva (Obinutuzumab), Fludarabine, Cyclophosphamide
35804589|T121|HDMP-R
35804589|T121|High Dose, MethylPrednisolone and Rituximab
35804589|T121|High Dose, MethylPrednisolone, Rituximab
35804590|T121|Idelalisib and Rituximab
35804590|T121|IdelaR
35804591|T121|Lenalidomide and Rituximab (R2)
35804591|T121|R<sup>2</sup>
35804591|T121|Rituximab and Revlimid (Lenalidomide)
35804591|T121|LR
35804592|T121|O-FC
35804592|T121|Ofatumumab, Fludarabine, Cyclophosphamide
35804593|T121|PCO
35804593|T121|Pentostatin, Cyclophosphamide, Ofatumumab
35804594|T121|Ofatumumab monotherapy
35804595|T121|PCR
35804595|T121|Pentostatin, Cyclophosphamide, Rituximab
35804595|T121|PER
35804595|T121|Pentostatin, Endoxan (Cyclophosphamide), Rituximab
35804596|T121|RCC
35804596|T121|Rituximab, Cladribine, Cyclophosphamide
35804597|T121|Non-curative first-line consolidation therapy
35804598|T121|Fludarabine monotherapy
35804598|T121|F
35804599|T121|CVP
35804599|T121|Cyclophosphamide, Vincristine, Prednisone
35804599|T121|Cyclophosphamide, Oncovin (Vincristine), Prednisone
35804599|T121|Vincristine, Cyclophosphamide, Prednisone
35804600|T121|R-FCM
35804600|T121|FCM-R
35804600|T121|Rituximab, Fludarabine, Cyclophosphamide, Mitoxantrone
35804600|T121|Fludarabine, Cyclophosphamide, Mitoxantrone, Rituximab
912006|T121|Ampicillin, Metronidazole, Bismuth
912007|T121|Antineoplastic monoclonal antibody
912008|T121|Anakinra
912009|T121|Ancestim
35804601|T121|Bendamustine and Rituximab (BR) and Ibrutinib
35804601|T121|BR and Ibrutinib
35804601|T121|Bendamustine, Rituximab, Ibrutinib
35804601|T121|IBR
35804601|T121|Ibrutinib, Bendamustine, Rituximab
35804602|T121|Bendamustine and Rituximab (BR) and Idelalisib
35804602|T121|BR and Idelalisib
35804602|T121|Bendamustine, Rituximab, Idelalisib
35804603|T121|Duvelisib monotherapy
35804604|T121|Idelalisib and Ofatumumab
35101853|T121|Andoprim
35804605|T121|Venetoclax and Rituximab
35804605|T121|VenR
35804606|T121|Acalabrutinib monotherapy
35804607|T121|Alemtuzumab and Rituximab
35804608|T121|Bendamustine and Ofatumumab
35804608|T121|BendOfa
35804609|T121|FluCam
35804610|T121|Fludarabine and Prednisone
35804611|T121|Ibrutinib and Ofatumumab
35804612|T121|Ibrutinib and Rituximab
35804613|T121|Idelalisib monotherapy
35804614|T121|Lenalidomide and Ofatumumab
35804615|T121|OFAR
35804615|T121|Oxaliplatin, Fludarabine, Ara-C (Cytarabine), Rituximab
35804616|T121|R-BAC
35804616|T121|Rituximab, Bendamustine, Ara-C (Cytarabine)
35804617|T121|Venetoclax monotherapy
35804618|T121|Non-curative subsequent-line consolidation therapy
35804619|T121|FC, then allo HSCT
35804619|T121|Fludarabine and Cyclophosphamide
35804620|T121|Fludarabine, Cyclophosphamide, ATG, then allo HSCT
35804621|T121|CAP
35804621|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Prednisone
35804622|T121|Chlorambucil monotherapy
35101852|T121|Anemul
35804623|T121|Chlorambucil and Prednisone
35804624|T121|Fludarabine and Rituximab (FR)
35804624|T121|FR
35804624|T121|Fludarabine and Rituximab
35804624|T121|Fludarabine, Rituximab
35804625|T121|Uracil mustard monotherapy
35101851|T121|Anitrim
35804626|T121|HDMP
35804626|T121|High Dose, MethylPrednisolone
912010|T121|Bendamustine and Dexamethasone
35804627|T121|Cytarabine and Interferon alfa-2b
35101850|T121|Anprim
912011|T121|Koselugo
35101849|T121|Ansentron
35101848|T121|Anset
35804628|T121|Hydroxyurea and Interferon alfa-2a
35804629|T121|Interferons
35101847|T121|Anti-CD79B antibody
911921|T121|CBM
35101846|T121|Antibac
35101845|T121|Anticoag
912012|T121|MET-mutated Non-small cell lung cancer
35804630|T121|Imatinib monotherapy, high dose
35804631|T121|Imatinib monotherapy, intermittent therapy
35804632|T121|Imatinib monotherapy, planned discontinuation
35804633|T121|Imatinib and LoDAC
35804633|T121|Imatinib and Low Dose Ara-C
35804634|T121|Imatinib and Interferon alfa
35804635|T121|Interferon alfa monotherapy
35804636|T121|Radotinib monotherapy
35804637|T121|BuCyTBI, then allo HSCT
35804637|T121|Busulfan, Cyclophosphamide, Total Body Irradiation
35804638|T121|Busulfan monotherapy
35101844|T121|Antrex
35101843|T121|Antrim
35101842|T121|Antrimox
912013|T121|Olaparib and Bevacizumab
912014|T121|Aripiprazole
35804639|T121|Interferon alfa-2b and DLI
35804639|T121|DLI
35804639|T121|Donor Lymphocyte Infusion
912015|T121|Atenolol
912016|T121|Pemazyre
912017|T121|INCB054828
912017|T121|Pemigatinib
35804640|T121|Omacetaxine monotherapy
35804641|T121| 2 Gy fractions x 27 fractions (total dose: 54 Gy), given 5 times per week, with boost to areas at high risk for malignant dissemination or that had inadequate resection margins of 2 Gy fractions x 6 fractions (boost dose: 12 Gy)
912018|T121|Pemigatinib monotherapy
35101841|T121|Apcetrim
35101840|T121|Aphtasolon
35101839|T121|Apidex
35804643|T121|Azacitidine and Lenalidomide
35804644|T121|Azacitidine and Vorinostat
35101838|T121|APO Sulfatrim
35804645|T121|Pletal
35804646|T121|Tagamet
35804647|T121|Cipro
35804648|T121|Abiplatin
35804649|T121|Axiplat
35804650|T121|Biocisplatinum
35804651|T121|Bioplatino
35804652|T121|Blastolem
35804653|T121|Briplatin
35804654|T121|Brisplatin
35804655|T121|C-Platin
35804656|T121|Ceplatin
35804657|T121|Ciplatan
35804658|T121|Ciplexal
35804659|T121|Cis-GRY
35804660|T121|Cismaplat
35804661|T121|Cispatin
35804662|T121|Cisplamerck
35804663|T121|Cisplan
35804664|T121|Cisplasol
35804665|T121|Cisplatex
35804666|T121|Cisplatine
35804667|T121|Cisplatino
35804668|T121|Cisplatyl
35804669|T121|Cisteen
35804670|T121|Citoplatino
35804671|T121|Cytoplatin
35804672|T121|Docistin
35804673|T121|Elvecis
35804674|T121|Fauldcispla
35804675|T121|Ifapla
35804676|T121|Kemoplat
35804677|T121|Lederplatin
35804678|T121|Metaplatin
35804679|T121|Neoplat
35804680|T121|Neoplatin
35804681|T121|Noveldexis
35804682|T121|Oncoplatin AQ
35804683|T121|Placis
35804684|T121|Platamin
35804685|T121|Platamine
35804686|T121|Platiblastin
35804687|T121|Platicis
35804688|T121|Platidiam
35804689|T121|Platikem
35804690|T121|Platil
35804691|T121|Platimit
35804692|T121|Platin
35804693|T121|Platinil
35804694|T121|Platino II Filaxis
35804695|T121|Platinol
35804696|T121|Platinox
35804697|T121|Platinoxan
35804698|T121|Platiran
35804699|T121|Platistil
35804700|T121|Platistin
35804701|T121|Platistine
35804702|T121|Platosin
35804703|T121|Randa
35804704|T121|Romcis
35804705|T121|Sicatem
35804706|T121|Sinplatin
35804707|T121|Sisplanil
35804708|T121|Tecnoplatin
35804709|T121|Tisplal
35804710|T121|Unistin
35804711|T121|Leustatin
35804712|T121|Litak
35804713|T121|Movectro
35804714|T121|Biaxin
35804715|T121|Clamist
35804716|T121|Dayhist
35804717|T121|Tavegil
35804718|T121|Tavist
35804719|T121|Clasteon
35804720|T121|Clastoban
35804721|T121|Climaclod
35804722|T121|Clodeosten
35804723|T121|Clodran
35804724|T121|Clodron
35804725|T121|Clody
35804726|T121|Difosfonal
35804727|T121|Disdual
35804728|T121|Lodronat
35804729|T121|Loron
35804730|T121|Lytos
35804731|T121|Mebonat
35804732|T121|Moticlod
35804733|T121|Niklod
35804734|T121|Ossiten
35804735|T121|Ostac
35804736|T121|Osteonorm
35804737|T121|Osteostab
35804738|T121|Sindronat
35804642|T121|Clolar
35804739|T121|Evoltra
35804740|T121|Evorabin
35804741|T121|Bio-Clopi
35804742|T121|Ceruvin
35804743|T121|Clop-75
35804744|T121|Clopalvix
35804745|T121|Clopicard
35804746|T121|Clopidro
35804747|T121|Clopinam
35804748|T121|Deviplat
35804749|T121|Lopigrol
35804750|T121|Plagril
35804751|T121|Plavix
35804752|T121|Stroka
35804753|T121|Cotellic
35101837|T121|APO-Bactotrim
912019|T121|Qinlock
35101836|T121|Apodrolen
35804754|T121|Colorectal cancer surgery
35804755|T121|CapeOx
35804755|T121|XELOX
35804755|T121|Capecitabine and Oxaliplatin
35804755|T121|XELoda (Capecitabine) and OXaliplatin
35804755|T121|CAPOX
35804755|T121|CAPecitabine and OXaliplatin
35804755|T121|CapeOX
35804755|T121|COX
35804755|T121|Capecitabine and OXaliplatin
35804755|T121|XELoda and OXaliplatin
35804755|T121|Capecitabine, OXaliplatin
35804755|T121|XELoda (Capecitabine), OXaliplatin
912020|T121|Retevmo
35101835|T121|Apotrinelax
912021|T121|DCC-2618
912021|T121|Ripretinib
912022|T121|Azacitidine IV monotherapy
912023|T121|Azacitidine oral monotherapy
912024|T121|Sacituzumab govitecan monotherapy
912025|T121|Azathioprine
912026|T121|LOXO-292
912026|T121|Selpercatinib
35101834|T121|Aptrim
35804756|T121|FLOX
35804756|T121|Fluorouracil, Leucovorin, OXaliplatin
35804757|T121|FOLFOX4
35804757|T121|FOLinic acid, Fluorouracil, OXaliplatin
35804757|T121|FOLinic acid, Fluorouracil, OXaliplatin 4
35804758|T121|mFOLFOX6
35804758|T121|modified FOLinic acid, Fluorouracil, OXaliplatin
35804758|T121|OxMdG
35804758|T121|Oxaliplatin Modified de Gramont
35804758|T121|FOLinic acid, Fluorouracil, OXaliplatin
912027|T121|MALT lymphoma
35804759|T121|Tegafur, Uracil, Folinic acid
35804759|T121|UFT + LV
35804759|T121|UFT (Tegafur and uracil) and LeucoVorin (Folinic acid)
35804760|T121|Metastasectomy
35804761|T121|FOLFIRI
35804761|T121|FOLinic acid, Fluorouracil, IRInotecan
35804761|T121|FUFIRI
35804761|T121|5-FU (Fluorouracil), Folinic acid, IRInotecan
35804761|T121|IF
35804761|T121|Irinotecan and 5-Fluorouracil
912028|T121|Tabrecta
35101833|T121|Aratran
35804762|T121|Surgery
35804763|T121|Hepatic arterial chemotherapy
35804764|T121|Intraperitoneal 5-FU
35804765|T121|Intraperitoneal hyperthermic mitomycin
912029|T121|Cytoreductive surgery
912030|T121|Trodelvy
912031|T121|Ixabepilone and Bevacizumab
912032|T121|Tukysa
35804766|T121|CapeOx and Bevacizumab
35804766|T121|CapeOX and Bevacizumab
35804766|T121|CAPOX-B
35804766|T121|XELOX and Bevacizumab
35804766|T121|Capecitabine, OXaliplatin, Bevacizumab
35804766|T121|CAPecitabine, OXaliplatin, Bevacizumab
35804766|T121|XELoda, OXaliplatin, Bevacizumab
912033|T121|ASTX727
912033|T121|Decitabine and cedazuridine
912034|T121|Decitabine and cedazuridine monotherapy
35804767|T121|CAPIRI
35804767|T121|CapeIRI
35804767|T121|XELIRI
35804767|T121|Capecitabine and IRInotecan
35804767|T121|CAPecitabine and IRInotecan
35804767|T121|XELox (Capecitabine) and IRInotecan
35804767|T121|mXELIRI
35804767|T121|modified XELox (Capecitabine) and IRInotecan
35804767|T121|XI
35804767|T121|Xeloda (Capecitabine) and Irinotecan
35804768|T121|CAPIRI-Bev
35804768|T121|XELIRI-Bev
35804768|T121|CAPecitabine, IRInotecan, Bevacizumab
35804768|T121|XELoda (Capecitabine), IRInotecan, Bevacizumab
35804768|T121|mXELIRI and Bevacizumab
35804768|T121|modified XELox (Capecitabine), IRInotecan, Bevacizumab
35804769|T121|Fluorouracil monotherapy
35101832|T121|Arcodexan
912035|T121|Bismuth subcitrate
912036|T121|Bismuth subsalicylate
912037|T121|E-CMF
912037|T121|Epirubicin followed by Cyclophosphamide, Methotrexate, Fluorouracil
35101831|T121|Arefarin
35101830|T121|Arendal
912038|T121|MFT
912039|T121|FEC-D
912039|T121|Fluorouracil, Epirubicin, Cyclophosphamide followed by Docetaxel
35804770|T121|FOLFIRI and Bevacizumab
35804770|T121|FOLinic acid, Fluorouracil, IRInotecan, Bevacizumab
35804771|T121|FOLFIRINOX
35804771|T121|FOLFOXIRI
35804771|T121|FOLinic acid, Fluorouracil, IRINotecan, OXaliplatin
35804771|T121|FOLinic acid, Fluorouracil, OXaliplatin, IRInotecan
35804771|T121|FFX
35804771|T121|Folinic acid, Fluorouracil, Irinotecan, Oxaliplatin
35804772|T121|FOLFIRINOX and Bevacizumab (L-Leucovorin)
35804772|T121|FOLFOXIRI and Bevacizumab
35804772|T121|L-FOLinic acid, Fluorouracil, IRINotecan, OXaliplatin, Bevacizumab
35804772|T121|L-FOLinic acid, Fluorouracil, OXaliplatin, IRInotecan, Bevacizumab
35804773|T121|FOLFOX2
35804773|T121|FOLinic acid, Fluorouracil, OXaliplatin
35101829|T121|Armol
912040|T121|Kitent
912041|T121|SHR-1210
912041|T121|HR-301210
912041|T121|Camrelizumab
35804774|T121|FOLFOX 7/sLV5FU2
35804774|T121|FOLinic acid, Fluorouracil, OXaliplatin alternating with simplified LeucoVorin, 5-FU, 2-weekly (every 2 weeks)
35804775|T121|mFOLFOX7
35804775|T121|modified FOLinic acid, Fluorouracil, OXaliplatin
35804776|T121|FOLFOX4 and Bevacizumab
35804776|T121|FOLFOX-B
35804776|T121|FOLinic acid, Fluorouracil, OXaliplatin, Bevacizumab
35804777|T121|mFOLFOX6-B
35804777|T121|FOLinic acid, Fluorouracil, OXaliplatin, Bevacizumab
35804777|T121|modified FOLinic acid, Fluorouracil, OXaliplatin, Bevacizumab
35804777|T121|FOLFOX-B
35804778|T121|IFL
35804778|T121|mIFL
35804778|T121|Irinotecan, Fluorouracil, Leucovorin (Folinic acid)
35804778|T121|modified Irinotecan, Fluorouracil, Leucovorin (Folinic acid)
912042|T121|Lenalidomide and Tafasitamab
35804779|T121|IFL and Bevacizumab
35804779|T121|mIFL and Bevacizumab
35804779|T121|Irinotecan, Fluorouracil, Leucovorin (Folinic acid), Bevacizumab
35804779|T121|modified Irinotecan, Fluorouracil, Leucovorin (Folinic acid), Bevacizumab
35804780|T121|IRIS and Bevacizumab
35804780|T121|IRInotecan, S-1, Bevacizumab
35804781|T121|IROX
35804781|T121|IRinotecan and OXaliplatin
35804782|T121|Nordic FLOX
35804782|T121|Fluorouracil, Leucovorin, OXaliplatin
35804783|T121|OXAFAFU
35804783|T121|OXAliplatin, Folinic Acid (Leucovorin), 5-FU (Fluorouracil)
35804784|T121|SOX
35804784|T121|S-1, OXaliplatin
35804784|T121|S-1 and OXaliplatin
912043|T121|Lucisun
35804785|T121|Non-curative second-line therapy
35101828|T121|Arond
35804786|T121|FOLFIRI and Ramucirumab
35804786|T121|FOLinic acid, Fluorouracil, IRInotecan and Ramucirumab
35804787|T121|FOLFIRI and Ziv-aflibercept
35804787|T121|FOLinic acid, Fluorouracil, IRInotecan, Ziv-aflibercept
912044|T121|Gavreto
35804788|T121|Non-curative third-line therapy
35804789|T121|Trifluridine and tipiracil monotherapy
35804790|T121|mFOLFOX6 and Cetuximab
35804790|T121|modified FOLinic acid, Fluorouracil, OXaliplatin, Cetuximab
35804790|T121|FOLFOX-C
35804790|T121|FOLinic acid, Fluorouracil, OXaliplatin, Cetuximab
42542272|T121|RAS wild-type Colorectal cancer
35804791|T121|CapeOx and Panitumumab
35804791|T121|Capecitabine, Oxaliplatin, Panitumumab
35804792|T121|FOLFIRI and Cetuximab
35804792|T121|FOLinic acid, Fluorouracil, IRInotecan, Cetuximab
35804793|T121|FOLFOX4 and Cetuximab
35804793|T121|FOLinic acid, Fluorouracil, OXaliplatin, Cetuximab
35804794|T121|FOLFOX4 and Panitumumab
35804794|T121|FOLinic acid, Fluorouracil, OXaliplatin, Panitumumab
35804795|T121|Cetuximab monotherapy
35804796|T121|mFOLFOXIRI and Cetuximab (L-Leucovorin)
35804796|T121|mFOLFOXIRI and Cetuximab
35804796|T121|modified L-FOLinic acid, Fluorouracil, OXaliplatin, IRInotecan, Cetuximab
35804797|T121|FOLFIRI and Panitumumab
35804797|T121|FOLinic acid, Fluorouracil, IRInotecan, Panitumumab
35804798|T121|Irinotecan and Cetuximab
35804799|T121| 2.0 Gy fractions given 5 times per week (total dose: 66-70 Gy)
912045|T121|Monjuvi
912046|T121|PGT
912047|T121|PGV
912048|T121|Clarithromycin, Metronidzole, PPI
35804800|T121|Panitumumab monotherapy
35804801|T121|Edrecolomab monotherapy
35804802|T121|Fluorouracil and Levamisole
912049|T121|Clarithromycin, Tetracycline, PPI, Bismuth
35804803|T121|FULV and Levamisole
35804803|T121|5-FU, LeucoVorin (Folinic acid), Levamisole
35804804|T121|MOF
35804804|T121|MeCCNU (Semustine), Oncovin (Vincristine), Fluorouracil
35804805|T121|Fluorouracil and Methotrexate (MF)
35804805|T121|Methotrexate and 5-Fluorouracil
35804806|T121|Fluorouracil and Mitomycin
35804807|T121|Fluorouracil and Semustine
35804808|T121|FOLFOX chronotherapy
35804808|T121|FOLinic acid, Fluorouracil, OXaliplatin
35804809|T121|Aliqopa
35804810|T121|Xalkori
35804811|T121|Belinostat monotherapy
35804812|T121|Bexarotene monotherapy
35804813|T121|Bexarotene and Pralatrexate
35804814|T121|Denileukin diftitox monotherapy
35804815|T121|Mogamulizumab monotherapy
35804816|T121|Pralatrexate monotherapy
35804817|T121|Romidepsin monotherapy
35804818|T121|Bleomycin and Cisplatin
35804819|T121|Cisplatin and Doxorubicin
35804819|T121|CD
35804819|T121|AP
35804819|T121|Adriamycin (Doxorubicin) and Platinol (Cisplatin)
35804819|T121|PLADO
35804819|T121|PLAtinol (Cisplatin) and DOxorubicin
35804820|T121|Sonidegib monotherapy
35804821|T121|Vismodegib monotherapy
35101827|T121|Ascotran
35804822|T121|Cemiplimab monotherapy
35804823|T121|Cisplatin, Interferon alfa-2a, Isotretinoin
35804824|T121|Berubigen
35804825|T121|CaloMist
35804826|T121|Cobavite
35804827|T121|Ener-B
35804828|T121|Nascobal
35804829|T121|Twelve Resin-K
35804830|T121|Alkyloxan
35804831|T121|Biodoxan
35804832|T121|Carloxan
35804833|T121|Ciclofosfamida
35804834|T121|Ciclokebir
35804835|T121|Cicloxal
35804836|T121|Clafen
35804837|T121|Claphene
35804838|T121|Cyclam
35804839|T121|Cycloblastin
35804840|T121|Cycloblastine
35804841|T121|CYCLO-cell
35804842|T121|Cycloferon
35804843|T121|Cyclomide
35804844|T121|Cyclophar
35804845|T121|Cyclophospham
35804846|T121|Cyclophosphamid
35804847|T121|Cyclophosphane
35804848|T121|Cyclostin
35804849|T121|Cyclostine
35804850|T121|Cyclotox
35804851|T121|Cycloxan
35804852|T121|Cycram
35804853|T121|Cydoxan
35804854|T121|Cyklofosfamid
35804855|T121|Cyphos
35804856|T121|Cytophosphan
35804857|T121|Cytoxan
35804858|T121|Cytoxan Lyophilized
35804859|T121|Endoxan
35804860|T121|Endoxan-N
35804861|T121|Endoxana
35804862|T121|Enduxan
35804863|T121|Formitex
35804864|T121|Fosfaseron
35804865|T121|Genoxal
35804866|T121|Genuxal
35804867|T121|Hidrofosmin
35804868|T121|Ledoxan
35804869|T121|Ledoxina
35804870|T121|Mitoxan
35804871|T121|Neophos
35804872|T121|Neosar
35804873|T121|Oncomide
35804874|T121|Oncophos
35804875|T121|Procytox
35804876|T121|Revimmune
35804877|T121|Sendoxan
35804878|T121|Siklofos
35804879|T121|Syklofosfamid
35804880|T121|Tymtran
35804881|T121|Zuviphos
35804882|T121|Zycram
35804883|T121|Zytoxan
35804884|T121|Gengraf
35804885|T121|Neoral
35804886|T121|Sandimmune
35804887|T121|Alcysten
35804888|T121|Alexan
35804889|T121|ARA
35804890|T121|Arabine
35804891|T121|Arabitin
35804892|T121|Aracitin
35804893|T121|Aracytin
35804894|T121|Aracytine
35804895|T121|Citagenin
35804896|T121|Citaloxan
35804897|T121|Citarabin
35804898|T121|Citarabina
35804899|T121|Citarabins
35804900|T121|Citarax
35804901|T121|Cylocide
35804902|T121|Cytarabin
35804903|T121|Cytarabins
35804904|T121|Cytarabinum
35804905|T121|Cytarbel
35804906|T121|Cytarine
35804907|T121|Cytosar
35804908|T121|Cytosar-U
35804909|T121|Cytrosar
35804910|T121|Depocyt
35804911|T121|Depocyte
35804912|T121|Erbabin
35804913|T121|Erpalfa
35804914|T121|Fauldcita
35804915|T121|Groven
35804916|T121|Ifarab
35804917|T121|Iretin
35804918|T121|Laracit
35804919|T121|Medsara
35804920|T121|Novutrax
35804921|T121|Remcyta
35804922|T121|Starasid
35804923|T121|Tabin
35804924|T121|Tabine
35804925|T121|Udicil
35804926|T121|Vyxeos
35804927|T121|Pradax
35804928|T121|Pradaxa
35804929|T121|Prazaxa
35804930|T121|Tafinlar
35804931|T121|Bazipar
35804932|T121|Cedcozine
35804933|T121|Dacarba
35804934|T121|Dacarex
35804935|T121|Dacin
35804936|T121|Dacmed
35804937|T121|Darbazine
35804938|T121|Dazine
35804939|T121|Decarb
35804940|T121|Oncodac
35804941|T121|Zydac
35804942|T121|Vizimpro
35804943|T121|Cosmegen
35804944|T121|Dacmozen
35804945|T121|Lyovac
35804946|T121|Daltepan
35804947|T121|Daltepin
35804948|T121|Fluzepamin
35804949|T121|Fragmin
35804950|T121|Fragmine
35804951|T121|Fragminject
35804952|T121|Fresubaru
35804953|T121|Hepachron
35804954|T121|Hepagumin
35804955|T121|Ligofragmin
35804956|T121|Low Liquemin
35804957|T121|Resolmin
35804958|T121|Orgaran
35804959|T121|Danatrol
35804960|T121|Danocrine
35804961|T121|Danodiol
35804962|T121|Danogen
35804963|T121|Drane
35804964|T121|Ladogal
35804965|T121|Novaprin
35804966|T121|Aczone
35804967|T121|Darzalex
35804968|T121|HuMax-CD38
35804969|T121|Actorise
35804970|T121|Aranesp
35804971|T121|Bionesp
35804972|T121|Cresp
35804973|T121|Darbetin
35804974|T121|Darbex
35804975|T121|Derise
35804976|T121|Kabidarba
35804977|T121|Nesp
35804978|T121|Nespo
35804979|T121|Sprycel
35804980|T121|Cerubidin
35804981|T121|Cerubidine
35804982|T121|D-Blastin
35804983|T121|Daunoblastin
35804984|T121|Daunoblastina
35804985|T121|Daunocin
35804986|T121|Daunomicina
35804987|T121|Daunorubicine
35804988|T121|Daurocina
35804989|T121|Maxidauno
35804990|T121|Ondena
35804991|T121|Rubidomycin
35804992|T121|Rubilem
35804993|T121|Rubomycin
35804994|T121|Runabicon
35804995|T121|DaunoXome
35804996|T121|Dacogen
35804997|T121|Decima
35804998|T121|Decita
35804999|T121|Decitafect
35805000|T121|Decitas
35805001|T121|Decitex
35805002|T121|Natdecita
35805003|T121|Exjade
35805004|T121|Jadenu
35805005|T121|Ferriprox
35805006|T121|Desferal
35805007|T121|Defitelio
35805008|T121|Firmagon
35805009|T121|Ontak
35805010|T121|Prolia
35805011|T121|Xgeva
35805012|T121|DDAVP
35805013|T121|DesmoMelt
35805014|T121|Desmotabs
35805015|T121|Desonap
35805016|T121|Minirin
35805017|T121|Stimate
35805018|T121|Dexam
35805019|T121|Oramin
35805020|T121|Polaramine
35805021|T121|Topmine
35805022|T121|Cardioxane
35805023|T121|Cyrdanax
35805024|T121|Savene
35805025|T121|Totect
35805026|T121|Zinecard
35805027|T121|R-ACVBP
35805027|T121|ACVBP-R
35805027|T121|Rituximab, Adriamycin (Doxorubicin), Cyclophosphamide, Vindesine, Bleomycin, Prednisone
35805027|T121|Adriamycin (Doxorubicin), Cyclophosphamide, Vindesine, Bleomycin, Prednisone, Rituximab
35805028|T121|R-CHOP
35805028|T121|R-CHOP-21
35805028|T121|CHOP-R
35805028|T121|RCHOP
35805028|T121|CHOPR
35805028|T121|Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone
35805028|T121|Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone given every 21 days
35805028|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone, Rituximab
35805028|T121|Rituximab, Cyclophosphamide, Hydroxydaunorubicin, Oncovin, Prednisone
35805028|T121|Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
35805028|T121|Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone every 21 days
35805029|T121|Orchiectomy
35805030|T121|Ibritumomab tiuxetan protocol
35101826|T121|Asmacortone
35805031|T121|R-CHOP-14
35805031|T121|Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone every 14 days
35805033|T121|R-MegaCHOP-14
35805033|T121|"Rituximab, ""Mega"" (high-dose) Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne every 14 days"
35805034|T121|R-miniCEOP
35805034|T121|Rituximab, mini, Cyclophosphamide, Epirubicin, O?? (vinblastine), Prednisone
35101825|T121|Asovorin
35805035|T121|Helicobacter pylori eradication therapy
35805036|T121|O-miniCHOP
35805036|T121|Ofatumumab, reduced-dose (<b>mini</b>) Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
35805037|T121|R-BL
35805037|T121|Rituximab, Bendamustine, Lenalidomide
35805037|T121|R2B
35805037|T121|Revlimid (Lenalidomide), Rituximab, Bendamustine
35805038|T121|R-CDOP
35805038|T121|DRCOP
35805038|T121|Rituximab, Cyclophosphamide, Doxil (Pegylated liposomal doxorubicin), Oncovin (Vincristine), Prednisone
35805038|T121|Doxil (Pegylated liposomal doxorubicin), Rituximab, Cyclophosphamide, Oncovin (Vincristine), Prednisone
35805038|T121|DR-COP
35805038|T121|Doxil (pegylated liposomal doxorubicin), Rituximab, Cyclophosphamide, Oncovin, Prednisone
35101824|T121|Aspen
35101823|T121|Aspirin and Warfarin
35805039|T121|R-CEOP90 (Epirubicin, Prednisolone)
35805039|T121|Rituximab, Cyclophosphamide, Epirubicin (90 mg/m<sup>2</sup> dosing), Oncovin (Vincristine), Prednisolone
35805032|T121|R-CEOP (Etoposide)
35805032|T121|R-CEOP
35805032|T121|Rituximab, Cyclophosphamide, Etoposide, Oncovin (Vincristine), Prednisone
35805040|T121|R-CHMP
35805040|T121|Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Marqibo (Vincristine liposomal), Prednisone
35805041|T121|R-GCVP
35805041|T121|Rituximab, Gemcitabine, Cyclophosphamide, Vincristine, Prednisolone
35805042|T121|R-MegaCHOP
35805042|T121|Rituximab, Mega, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
35805043|T121|R-IFE
35805043|T121|REI
35805043|T121|Rituximab, IFosfamide, Etoposide
35805043|T121|Rituximab, Etoposide, Ifosfamide
35805044|T121|R-miniCHOP
35805044|T121|Rituximab, reduced-dose (<b>mini</b>) Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
35805045|T121|R2-CHOP
35805045|T121|LR-CHOP-21
35805045|T121|Rituximab, Revlimid (Lenalidomide), Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone
35805045|T121|Lenalidomide, Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone given every 21 days
35805046|T121|Low molecular weight heparins
35805047|T121|CBV, then auto HSCT
35805048|T121|CBVM
35805049|T121|ACE
35805049|T121|Adriamycin (Doxorubicin), Cyclophosphamide, Etoposide
35805049|T121|AVE
35805049|T121|CAE
35805049|T121|Adriamycin (Doxorubicin), Vepesid (Etoposide), Endoxan (Cyclophosphamide)
35805049|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Etoposide
35805050|T121|ACVBP
35805050|T121|Adriamycin (Doxorubicin), Cyclophosphamide, Vindesine, Bleomycin, Prednisone
35805051|T121|Z-BEAM, then auto HSCT
35805052|T121|O-DHAP
35805052|T121|Ofatumumab, Dexamethasone, High-dose Ara-C (Cytarabine), Platinol (Cisplatin)
35101822|T121|Assepium
35805053|T121|O-ICE
35805053|T121|Ofatumumab, Ifosfamide, Carboplatin, Etoposide
35805054|T121|R-DexaBEAM
35805054|T121|Rituximab, Dexamethasone, BiCNU (Carmustine), Etoposide, Ara-C (Cytarabine), Melphalan
35805055|T121|R-BEAM, then auto HSCT
35805056|T121|R-TBI/Cy, then auto HSCT
35805057|T121|R-DHAOx
35805057|T121|ROAD
35805057|T121|Rituximab, Dexamethasone, High-dose Ara-C (Cytarabine), Oxaliplatin
35805057|T121|Rituximab, Oxaliplatin, Ara-C (Cytarabine), Dexamethasone
35805058|T121|R-DHAP
35805058|T121|Rituximab, Dexamethasone, High-dose Ara-C (Cytarabine), Platinol (Cisplatin)
35805059|T121|R-DHAP/R-VIM
35805059|T121|Rituximab, Dexamethasone, High-dose Ara-C (Cytarabine), Platinol (Cisplatin) alternating with Rituximab, VP-16 (Etoposide), Ifosfamide, Methotrexate
35805060|T121|R-EPOCH
35805060|T121|Rituximab, Etoposide, Prednisone, Oncovin (Vincristine), Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin)
35805061|T121|R-ESHAP
35805061|T121|Rituximab, Etoposide, Solumedrol (Methylprednisolone) High-dose Ara-C (Cytarabine), Platinol (Cisplatin)
35805062|T121|R-GDP
35805062|T121|Rituximab, Gemcitabine, Dexamethasone, Platinol (Cisplatin)
35805063|T121|R-ICE
35805063|T121|ICE-R
35805063|T121|Rituximab, Ifosfamide, Carboplatin, Etoposide
35805063|T121|Ifosfamide, Carboplatin, Etoposide, Rituximab
35805064|T121|RICER
35805064|T121|Rituximab, Ifosfamide, Carboplatin, Etoposide, Revlimid (Lenalidomide)
35805065|T121|R-NIMP
35805065|T121|Rituximab, Navelbine (Vinorelbine), Ifosfamide, Mitoxantrone, Prednisone
35805066|T121|BEAC, then auto HSCT
35805067|T121|BEAM, then allo HSCT
35805067|T121|BiCNU (Carmustine), Etoposide, Ara-C (Cytarabine), Melphalan
35805068|T121|BeEAM, then auto HSCT
35805069|T121|Cyclophosphamide and TBI, then auto HSCT
35805070|T121|FEAM, then auto HSCT
35805071|T121|Fludarabine, Busulfan, ATG, Ibritumomab tiuxetan, then allo HSCT
35805072|T121|LEED, then auto HSCT
912050|T121|TCHL (Docetaxel)
35805073|T121|Maintenance after salvage therapy
912051|T121|TCL (Docetaxel)
35805074|T121|Axicabtagene ciloleucel monotherapy
912052|T121|Cytotoxic chemotherapeutic
35805075|T121|Everolimus monotherapy
35805076|T121|Everolimus and Rituximab
35805077|T121|GVD
35805077|T121|Gemcitabine, Vinorelbine, Doxil (Pegylated liposomal doxorubicin)
35101821|T121|Athrombin-K
35805078|T121|Oxaliplatin monotherapy
35805079|T121|Panobinostat and Rituximab
35805080|T121|Pixantrone monotherapy
35101820|T121|Atomexin
35805081|T121|R-CVEP
35805081|T121|Rituximab, Cyclophosphamide, Vorinostat, Etoposide, Prednisone
35101819|T121|Atossa
35805082|T121|R-GemOx
35805082|T121|Rituximab, Gemcitabine, Oxaliplatin
35805082|T121|GEMOX-R
35805082|T121|GEMcitabine, OXaliplatin, Rituximab
35805083|T121|R-INO
35805083|T121|Rituximab, INOtuzumab ozogamicin
35805084|T121|TTR
35805084|T121|Taxol (Paclitaxel), Topotecan, Rituximab
35805085|T121|ABP
35805085|T121|Adriamycin (Doxorubicin), Bleomycin, Prednisone
35805086|T121|ACOMLA
35805086|T121|Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Methotrexate, Leucovorin (Folinic acid), Ara-C (Cytarabine)
35805087|T121|BCOP
35805087|T121|BCNU (Carmustine), Cyclophosphamide, Oncovin (Vincristine), Prednisone
35805088|T121|CAP-BOP
35805088|T121|COP-BLAM
35805088|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Procarbazine, Bleomycin, Oncovin (Vincristine), Prednisone
35805088|T121|Cyclophosphamide, Oncovin (Vincristine), Prednisone, BLeomycin, Adriamycin (Doxorubicin), Matulane (Procarbazine),
35805089|T121|CCOP
35805089|T121|Cyclophosphamide, Caelyx (Pegylated liposomal doxorubicin), Oncovin (Vincristine), Prednisone
35805090|T121|CEEP
35805090|T121|Cyclophosphamide, Epirubicin, Eldesine (Vindesine), Prednisone
35805091|T121|CEOP
35805091|T121|Cyclophosphamide, Epirubicin, Oncovin (Vincristine), Prednisone
35805092|T121|CHOP Modified
35805092|T121|mCHOP
35805092|T121|modified Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone
35805093|T121|CHOP-BCG
35805093|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone, Bacillus Calmette-Guerin
35805094|T121|CHOP-B
35805094|T121|B-CHOP
35805094|T121|BACOP
35805094|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone, Bleomycin
35805094|T121|Bleomycin, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone
35805094|T121|Bleomycin, Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Prednisone
35805094|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne, Bleomycin
35805095|T121|C-MOPP
35805095|T121|COPP
35805095|T121|CyclophosphaMide, Oncovin (Vincristine), Procarbazine, Prednisone
35805095|T121|Cyclophosphamide, Oncovin (Vincristine), Procarbazine, Prednisone
35805096|T121|CNOP
35805096|T121|MCOP
35805096|T121|Cyclophosphamide, Novantrone (Mitoxantrone), Oncovin (Vincristine), Prednisone
35805096|T121|Mitoxantrone, Cyclophosphamide, Oncovin (Vincristine), Prednisone
35805097|T121|COP-Bleo
35805097|T121|Cyclophosphamide, Oncovin (Vincristine), Prednisone, Bleomycin
35101818|T121|Auxiloson
35805098|T121|DICEP
35805098|T121|Dose Intensive Cyclophosphamide, Etoposide, Platinol (Cisplatin)
35805099|T121|F-MACHOP
35805099|T121|Fluorouracil, Methotrexate, Ara-C (Cytarabine), Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
35101817|T121|Auxison
35101816|T121|Auxisone
35101815|T121|Avancort
35805100|T121|HOP
35805100|T121|Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone
35805100|T121|Adriamycin (Doxorubicin), Prednisone, Oncovin (Vincristine)
35805101|T121|LD-ACOP-B
35805101|T121|Low-Dose Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Prednisone, Bleomycin
35805102|T121|MACOP-B
35805102|T121|Methotrexate, Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Prednisone, Bleomycin
35101814|T121|Avlotrin
35805103|T121|m-BACOD
35805103|T121|methotrexate (moderate dose), Bleomycin, Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Dexamethasone
35805104|T121|m-BNCOD
35805104|T121|methotrexate (moderate dose), Bleomycin, Novantrone (Mitoxantrone), Cyclophosphamide, Oncovin (Vincristine), Dexamethasone
35805105|T121|P/DOCE
35805105|T121|Prednisone, Doxorubicin, Oncovin (Vincristine), Cyclophosphamide, Etoposide,
35805106|T121|PACEBOM
35805106|T121|Prednisolone, Adriamycin (Doxorubicin), Cyclophosphamide, Etoposide, Bleomycin, Oncovin (Vincristine), Methotrexate
35805107|T121|PEN
35805107|T121|Prednisone, Etoposide, Novantrone (Mitoxantrone)
35805108|T121|PMitCEBO
35805108|T121|Prednisolone, Mitoxantrone, Cyclophosphamide, Etoposide, Bleomycin, Oncovin (Vincristine)
35101813|T121|Axitinib and Pembrolizumab
42542273|T121|CAFVP
42542273|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Fluorouracil, Vincristine, Prednisone
35805109|T121|ProMACE-CytaBOM
35805109|T121|Prolix (Prednisone), Methotrexate, Adriamycin (Doxorubicin), Cyclophosphamide, Etoposide, Cytarabine, Bleomycin, Oncovin (Vincristine), Methotrexate
35805110|T121|ProMACE-MOPP
35805110|T121|Prolix (Prednisone), Methotrexate, Adriamycin (Doxorubicin), Cyclophosphamide, Etoposide, Mustargen (Mechlorethamine), Oncovin (Vincristine), Procarbazine, Prednisone
35805111|T121|VABE
35805111|T121|Vincristine, Adriamycin (Doxorubicin), Bleomycin, Etoposide, Prednisone
35805112|T121|VACOP-B
35805112|T121|P-VABEC
35805112|T121|Vepesid (Etoposide), Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Prednisone, Bleomycin
35805112|T121|Prednisone, Vincristine, Adriamycin (Doxorubicin), Bleomycin, Etoposide, Cyclophosphamide
35805113|T121|VCAP
35805113|T121|Vindesine, Cyclophosphamide, Adriamycin (Doxorubicin), Prednisone
35805114|T121|VEPA
35805114|T121|Vincristine, Endoxan (Cyclophosphamide), Prednisolone, Adriamycin (Doxorubicin)
35805115|T121|VNCOP-B
35805115|T121|Vepesid (Etoposide), Novantrone (Mitoxantrone), Cyclophosphamide, Oncovin (Vincristine), Prednisone, Bleomycin
35805116|T121|VR-CHOP
35805116|T121|RB-CHOP
35805116|T121|Velcade (Bortezomib), Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
35805116|T121|Rituximab, Bortezomib, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
35805116|T121|Velcade (Bortezomib) Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
35805117|T121|EPIC regimen
35805117|T121|Etoposide, Prednisolone, Ifosfamide, Carboplatin
35805118|T121|MINE
35805118|T121|Mesna, Ifosfamide, Novantrone (Mitoxantrone), Etoposide
35805119|T121|ESHAP
35805119|T121|Etoposide, Solumedrol (Methylprednisolone), High dose Ara-C (Cytarabine), Platinol (Cisplatin)
35805119|T121|Etoposide, Solumedrol (Methylprednisolone) High-dose Ara-C (Cytarabine), Platinol (Cisplatin)
35805120|T121|VIM
35805120|T121|Vepesid (Etoposide), Ifosfamide, Mitoxantrone
35805121|T121|VIPD
35805121|T121|DVIP
35805121|T121|VP-16 (Etoposide), Ifosfamide, Platinol (Cisplatin), Dexamethasone
35805121|T121|Dexamethasone, VP-16 (Etoposide), Ifosfamide, Platinol (Cisplatin)
35805122|T121|CEPP(B)
35805122|T121|Cyclophosphamide, Etoposide, Procarbazine, Prednisone, (optional) Bleomycin
35805123|T121|DICE
35805123|T121|Dexamethasone, Ifosfamide, Carboplatin, Etoposide
35805124|T121|EPOCH
35805124|T121|CHEOP
35805124|T121|Etoposide, Prednisone, Oncovin (Vincristine), Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin)
35805124|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Etoposide, Oncovin (Vincristine), Prednisone
35805125|T121|Etoposide, Ifosfamide, Methotrexate
35805125|T121|IMVP-16
35805125|T121|Ifosfamide, Methotrexate, VP-16 (Etoposide)
35805126|T121|ICE
35805126|T121|Ifosfamide, Carboplatin, Etoposide
35805127|T121|Unituxin
35805128|T121|Benadryl
35805129|T121|Persantine
35805130|T121|Asodocel
35805131|T121|Daxotel
35805132|T121|Docefrez
35805133|T121|Docegem
35805134|T121|Doceglob
35805135|T121|Docemax
35805136|T121|Docenat
35805137|T121|Docepar
35805138|T121|Docetax
35805139|T121|Docetec
35805140|T121|Docetere
35805141|T121|DoceXan
35805142|T121|Docshil
35805143|T121|Dolectran
35805144|T121|Doxel
35805145|T121|Doxetal
35805146|T121|Hentaxel
35805147|T121|Neocel
35805148|T121|Oncodocel
35805149|T121|Plustaxano
35805150|T121|Sibatere
35805151|T121|Taceedo
35805152|T121|Taxe-RTU
35805153|T121|Taxewell
35805154|T121|Taxotere
35805155|T121|Texot
35805156|T121|Trixotene
35805157|T121|Uvtere
35805158|T121|Colace
35805159|T121|Anzemet
35805160|T121|Motilium
35805161|T121|Didox
35805162|T121|Adriablastina
35805163|T121|Adriacept
35805164|T121|Adriacin
35805165|T121|Adriamycin
35805166|T121|Adriblastin
35805167|T121|Adriblastina
35805168|T121|Adriblastine
35805169|T121|Adricept
35805170|T121|Adricin
35805171|T121|Adrim
35805172|T121|Adrimedac
35805173|T121|Adrosal
35805174|T121|Antraciclin
35805175|T121|Biorrub
35805176|T121|Biorubina
35805177|T121|Cadria
35805178|T121|Carcinocin
35805179|T121|Cloridrato DE
35805180|T121|Doxorrubicina Colhidrol
35805181|T121|Deldoxin
35805182|T121|Dicladox
35805183|T121|Dobicin
35805184|T121|Dobixin
35805185|T121|Doxo
35805186|T121|Doxobin
35805187|T121|Doxo Cell
35805188|T121|Doxocris
35805189|T121|Doxokebir
35805190|T121|Doxolem
35805191|T121|Doxonolver
35805192|T121|Doxor
35805193|T121|Doxorrubicina
35805194|T121|Doxoruben
35805195|T121|Doxorubicina
35805196|T121|Doxorubicine
35805197|T121|Doxorubicinum
35805198|T121|Doxorubin
35805199|T121|Doxotec
35805200|T121|Doxtie
35805201|T121|Duxocin
35805202|T121|Evacet
35805203|T121|Farmiblastina
35805204|T121|Fauldoxo
35805205|T121|Flavicina
35805206|T121|Ifadox
35805207|T121|Kemodoxa
35805208|T121|Lipodox
35805209|T121|Lyphidox
35805210|T121|Myocet
35805211|T121|Nagun
35805212|T121|Neoxane
35805213|T121|Nuaze
35805214|T121|Oncodria
35805215|T121|Onkodox
35805216|T121|Onkostatil
35805217|T121|Pallagicin
35805218|T121|Ranxas
35805219|T121|Rastocin
35805220|T121|Ribodoxo
35805221|T121|Roxorin
35805222|T121|Rubex
35805223|T121|Varidoxo
35805224|T121|Zodox
35805225|T121|Marinol
35805226|T121|Imfinzi
35805227|T121|Avodart
35805228|T121|Copiktra
35805229|T121|Erlotinib monotherapy
42542274|T121|EGFR-mutated malignancy
35805230|T121|Ado-trastuzumab emtansine monotherapy
42542275|T121|ERBB2-mutated malignancy
42542276|T121|ERBB3-mutated malignancy
35805231|T121|Soliris
35805232|T121|Savaysa
35805233|T121|Panorex
35805234|T121|Empliciti
35805235|T121|Eltrom
35805236|T121|Promacta
35805237|T121|Revolade
35805238|T121|Hemlibra
35805239|T121|Idhifa
35805240|T121|Braftovi
35805241|T121|Endocrine ablation surgery
35805242|T121|Endometrial cancer surgery
35805243|T121|CIM
35805243|T121|Cisplatin, Ifosfamide, Mesna
35805244|T121|Whole abdominal radiation (WAI)
35805245|T121|Carboplatin and Pegylated liposomal doxorubicin
35805245|T121|CD
35805245|T121|PLDC
35805245|T121|Carboplatin and Doxil (Pegylated liposomal doxorubicin)
35805245|T121|Pegylated Liposomal Doxorubicin and Carboplatin
35805246|T121|Cisplatin, Doxorubicin, Paclitaxel
35805246|T121|TAP
35805246|T121|Taxol (Paclitaxel), Adriamycin (Doxorubicin), Platinol (Cisplatin)
35805247|T121|Dactinomycin monotherapy
35101812|T121|B Dexzol
35805248|T121|Ifosfamide and Paclitaxel
35805248|T121|PI
35805248|T121|Paclitaxel and Ifosfamide
35805248|T121|Paclitaxel, Ifosfamide
35805248|T121|TI
35805248|T121|Taxol (Paclitaxel) and Ifosfamide
35101811|T121|B.S.
35805249|T121|Medroxyprogesterone and Tamoxifen
35805250|T121|Megestrol and Tamoxifen
35805251|T121|Axoparin
35805252|T121|Cardinex
35805253|T121|Clexan
35805254|T121|Clexane
35805255|T121|Clotinex
35805256|T121|Cnoxane
35805257|T121|Cutenox
35805258|T121|Dutenox
35805259|T121|Enclex
35805260|T121|Enox
35805261|T121|Enxoaealth
35805262|T121|Enoxol
35805263|T121|Eparin
35805264|T121|Lmwx
35805265|T121|Lovenox
35805266|T121|Markparin
35805267|T121|Microparin
35805268|T121|Noxprin
35805269|T121|Pariparin
35805270|T121|Xaparin
35805271|T121|Xtandi
35805272|T121|Alrubicin
35805273|T121|Anthracin
35805274|T121|Binarin
35805275|T121|Bioepicyna
35805276|T121|Crisabon
35805277|T121|E.P.R Elvetium
35805278|T121|Ellence
35805279|T121|Epidoxo
35805280|T121|Epifil
35805281|T121|Epilem
35805282|T121|Epirubicine
35805283|T121|Epizin
35805284|T121|Epricin
35805285|T121|Eracin
35805286|T121|Famorubicin
35805287|T121|Farmorubicin
35805288|T121|Farmorubicina
35805289|T121|Farmorubicine
35805290|T121|Pharmorubicin
35805291|T121|Riboepi
35805292|T121|Rubifarm
35805293|T121|Retacrit
35805294|T121|Ceriton
35805295|T121|Dynepo
35805296|T121|Epoch
35805297|T121|Epofer
35805298|T121|Epogen
35805299|T121|Epogin
35805300|T121|Epoimmun
35805301|T121|Epomax
35805302|T121|Epopen
35805303|T121|Epox
35805304|T121|Epoyet
35805305|T121|Eprex
35805306|T121|Eritrelan
35805307|T121|Erypo
35805308|T121|Erythrostim
35805309|T121|Espo
35805310|T121|Globuren
35805311|T121|Hemapo
35805312|T121|Hemax
35805313|T121|LG Espogen
35805314|T121|Procrit
35805315|T121|Recormon
35805316|T121|Vepox
35805317|T121|Vintor
35805318|T121|Wepox
35805319|T121|Integrilin
35805320|T121|Balversa
35805321|T121|Cobimetinib monotherapy
35805322|T121|Sirolimus and Prednisone
35805323|T121|Halaven
35805324|T121|Erlocip
35805325|T121|Erlonat
35805326|T121|Melacyte
35805327|T121|Tarceva
35805328|T121|Cisplatin, Docetaxel, RT
35805328|T121|DC and RT
35805328|T121|Docetaxel, Cisplatin, Radiation Therapy
35805328|T121|DP and RT
35805328|T121|Docetaxel, Platinol (Cisplatin), Radiation Therapy
35805329|T121|Cisplatin and Etoposide (EP)
35805329|T121|PE
35805329|T121|EC
35805329|T121|Platinol (Cisplatin) and Etoposide
35805329|T121|Etoposide and Cisplatin
35805329|T121|Etoposide, Platinol (Cisplatin)
35805329|T121|Etoposide and Platinol (Cisplatin)
35805329|T121|Platinol (Cisplatin), Etoposide
35805330|T121|Esophageal cancer surgery
35805331|T121|Fluorouracil, Paclitaxel, RT
35805331|T121|Fluorouracil, Paclitaxel, Radiation Therapy
35805332|T121|Cisplatin, Irinotecan, RT
35805332|T121|Cisplatin, Irinotecan, Radiation Therapy
35101810|T121|BAC-Sulfitrin
35805333|T121|CLF
35805333|T121|PLF
35805333|T121|Cisplatin, Leucovorin (Folinic acid), Fluorouracil
35805333|T121|Platinol (Cisplatin), Leucovorin (Folinic acid), Fluorouracil
35805333|T121|FLP
35805333|T121|Cisplatin, Leucovorin, Fluorouracil
35805333|T121|Fluorouracil, Leucovorin, Platinol (Cisplatin)
35805334|T121|Cisplatin, Etoposide, RT
35805334|T121|EP and RT
35805334|T121|Etoposide, Platinol (Cisplatin), Radiation Therapy
35805334|T121|PE + RT
35805334|T121|Platinol (Cisplatin), Etoposide, Radiation Therapy
35805335|T121|Capecitabine and Cisplatin (CX)
35805335|T121|CX
35805335|T121|XP
35805335|T121|Cisplatin and Xeloda (Capecitabine)
35805335|T121|Xeloda (Capecitabine) and Platinol (Cisplatin)
35805335|T121|Cisplatin, Xeloda (Capecitabine)
35805335|T121|Xeloda (Capecitabine), Platinol (Cisplatin)
35805336|T121|Capecitabine, Cisplatin, RT
35805336|T121|CX and RT
35805336|T121|Cisplatin, Xeloda (Capecitabine), Radiation Therapy
35805337|T121|ECX
35805337|T121|Epirubicin, Cisplatin, Xeloda (Capecitabine)
35805337|T121|ECC
35805337|T121|Epirubicin, Cisplatin, Capecitabine
35805338|T121|EOF
35805338|T121|Epirubicin, Oxaliplatin, Fluorouracil
35805338|T121|Epirubicin, Oxaliplatin, Fluourouracil
35805339|T121|EOX
35805339|T121|EOC
35805339|T121|Epirubicin, Oxaliplatin, Xeloda (Capecitabine)
35805339|T121|Epirubicin, Oxaliplatin, Capecitabine
35805340|T121|FLEP
35805340|T121|Fluorouracil, Leucovorin, Etoposide, Platinol (Cisplatin)
35101809|T121|Bacfar
35805341|T121|FLOT
35805341|T121|Fluorouracil, Leucovorin, Oxaliplatin, Taxotere (Docetaxel)
35805342|T121|PCF
35805342|T121|Paclitaxel, Cisplatin, Fluorouracil
35805342|T121|PPF
35805342|T121|Paclitaxel, Platinol (Cisplatin), Fluorouracil
35805343|T121|Capecitabine, Carboplatin, Paclitaxel, RT
35805343|T121|Capecitabine, Carboplatin, Paclitaxel, Radiation Therapy
35805344|T121|Esophagectomy
35805345|T121|Capecitabine, Docetaxel, RT
35805345|T121|Capecitabine, Docetaxel, Radiation Therapy
35805346|T121|Capecitabine, Docetaxel, Oxaliplatin, RT
35805346|T121|Capecitabine, Docetaxel, Oxaliplatin, Radiation Therapy
35805347|T121|Capecitabine, Oxaliplatin, RT
35805347|T121|Capecitabine, Oxaliplatin, Radiation Therapy
35805348|T121|Capecitabine, Paclitaxel, RT
35805348|T121|Capecitabine, Paclitaxel, Radiation Therapy
35805349|T121|Carboplatin, Fluorouracil, RT
35805349|T121|Carboplatin, Fluorouracil, Radiation Therapy
35805350|T121|Carboplatin and Paclitaxel (CP) and RT
35805350|T121|CP and RT
35805350|T121|"<table class=""wikitable"" style=""color:black; background-color:#42f584"">"
35805350|T121|Carboplatin, Paclitaxel, Radiation Therapy
35805350|T121|Carboplatin, Paclitaxel, RT
35805350|T121|PC and RT
35805350|T121|Paclitaxel, Carboplatin, Radiation Therapy
912053|T121|Neutrexin
35101808|T121|Bacidal
35805351|T121|Cisplatin, Vinorelbine, RT
35805351|T121|Cisplatin, Vinorelbine, Radiation Therapy
35805352|T121|Docetaxel, Fluorouracil, RT
35805352|T121|Docetaxel, Fluorouracil, Radiation Therapy
35805353|T121|Fluorouracil, Oxaliplatin, RT
35805353|T121|Fluorouracil, Oxaliplatin, Radiation Therapy
35101807|T121|Bacin
35101806|T121|Bacitran
35101805|T121|Bacmetrin
35101804|T121|Bacoprim
35101803|T121|Bacotrin
912054|T121|Onureg
35101802|T121|Bacprotin
35101801|T121|Bacris
35805354|T121|FOLFOX4 and RT
35805354|T121|FOLinic acid, Fluorouracil, OXaliplatin, Radiation Therapy
35805355|T121|5-FU and Leucovorin, then 5-FU, Leucovorin, RT, then 5-FU and Leucovorin
35805356|T121|ECF/5-FU and RT
35805356|T121|Epirubicin, Cisplatin, Fluorouracil alternating with 5-FluoroUracil and Radiation Therapy
35101800|T121|Bacsulfaprin
35805357|T121|Apatinib monotherapy
35101799|T121|Bacsultrim
35101798|T121|Bactar
35101797|T121|Bactazol
35101796|T121|Bactekod
35101795|T121|Bactelan
35805358|T121|Carboplatin, Docetaxel, Fluorouracil
35101794|T121|Bacteracin
35101793|T121|Bacterial
35101792|T121|Bacteric
912055|T121|Pixantrone and Rituximab
35805359|T121|Cisplatin and Fluorouracil (CF) and Cetuximab
35805359|T121|CF-C
35805359|T121|Cisplatin, Fluorouracil, Cetuximab
35805360|T121|Cisplatin and Fluorouracil (CF) and Trastuzumab
35805360|T121|CF and Trastuzumab
35805360|T121|Cisplatin, Fluorouracil, Trastuzumab
35805361|T121|LdCF
35805361|T121|Liposomal doxorubicin, Cisplatin, Fluorouracil
35101791|T121|Bacteriof.klebs PN
912056|T121|Danyelza
35101790|T121|Bacterol
35101789|T121|Bacticel
35101788|T121|Bactide
35101787|T121|Bactifor
35101786|T121|Bactigram
35101785|T121|Bactille-TS
35805362|T121|CX-C
35805363|T121|Capecitabine and Cisplatin (CX) and Trastuzumab
35805363|T121|CX and Trastuzumab
35805363|T121|Cisplatin, Xeloda (Capecitabine), Trastuzumab
35101784|T121|Bactipront
35101783|T121|Bactiseptol
912057|T121|TAK-385
912057|T121|Relugolix
35805364|T121|DCF
35805364|T121|Docetaxel, Cisplatin, Fluorouracil
35805364|T121|TCF
35805364|T121|Taxotere (Docetaxel), Cisplatin, Fluorouracil
35805364|T121|TPF
35805364|T121|Taxotere (Docetaxel), Platinol (Cisplatin), Fluorouracil
35101782|T121|Bactiver
912058|T121|Dara-CyBorD
912058|T121|D-VCd
912058|T121|Daratumumab and hyaluronidase, Cyclophosphamide, Bortezomib, Dexamethasone
912058|T121|Daratumumab and hyaluronidase, Velcade (Bortezomib), Cyclophosphamide, low-dose dexamethasone
35101781|T121|Bactoprim
35805365|T121|mDCF and Bevacizumab
35805365|T121|modified Docetaxel, Cisplatin, Fluorouracil and Bevacizumab
35805366|T121|Docetaxel and Irinotecan
35101780|T121|Bactoreduct
35805367|T121|DOF
35101779|T121|Bactosain
912059|T121|RET-positive Non-small cell lung cancer
35101778|T121|Bactostab
912060|T121|RET-positive Thyroid cancer
35101777|T121|Bactramin
912061|T121|Ripretinib monotherapy
35101776|T121|Bactricid
35101775|T121|Bactricida
35101774|T121|Bactricin
35101773|T121|Bactrilac
35101772|T121|Bactrim
35101771|T121|Bactrimel
35101770|T121|Bactrin
35805368|T121|Irinotecan liposomal monotherapy
35805369|T121|Irinotecan and Mitomycin
35101769|T121|Bactrisan
35101768|T121|Bactrium DS
35101767|T121|Bactrizole
35805370|T121|MCF
35805370|T121|Mitomycin, Cisplatin, Fluorouracil
35101766|T121|Bactron
35101765|T121|Bactronil
912062|T121|Selpercatinib monotherapy
35805371|T121|Paclitaxel and Ramucirumab
35101764|T121|Bactropin
35805372|T121|Ramucirumab monotherapy
35805373|T121|Anagrelide monotherapy
35805374|T121|Aspirin and Anagrelide
912063|T121|Sunitix
35805375|T121|Aspirin and Hydroxyurea
35805376|T121|Hydroxyurea monotherapy
35101763|T121|Bacxal
35805377|T121|Peginterferon alfa-2a monotherapy
35101762|T121|Baczin
35101761|T121|Baczole
35805380|T121|Emcyt
35805381|T121|Estracit
35805382|T121|Estram
35805383|T121|Estramin
35805384|T121|X-Trant
35805385|T121|Aside
35805386|T121|Beposid
35805387|T121|Bioposide
35805388|T121|Celltop
35805389|T121|Citodox
35805390|T121|Epocin
35805391|T121|Eposid
35805392|T121|Eposide
35805393|T121|Eposido
35805394|T121|Eposin
35805395|T121|Epsidox
35805396|T121|ETO
35805397|T121|Etocris
35805398|T121|Etomedac
35805399|T121|Etonolver
35805400|T121|Etopofos
35805401|T121|Etopophos
35805402|T121|Etopos
35805403|T121|Etoposid
35805404|T121|Etoposido
35805405|T121|Etopoxan
35805406|T121|Etopul
35805407|T121|Etosid
35805408|T121|Etosin
35805409|T121|Eunades CS
35805410|T121|Euvaxon
35805411|T121|Exitop
35805412|T121|Fytop
35805413|T121|Fytosid
35805414|T121|Labimion
35805415|T121|Lastet
35805416|T121|Lastet S
35805417|T121|Neoplaxol
35805418|T121|Nexvep
35805419|T121|Onkoposid
35805420|T121|Optasid
35805421|T121|Percas
35805422|T121|Posid
35805423|T121|Posidon
35805424|T121|Posyd
35805425|T121|Riboposid
35805426|T121|Sintopozid
35805427|T121|Toposar
35805428|T121|Toposide
35805429|T121|Toposin
35805430|T121|Topresid
35805431|T121|Tosuben
35805432|T121|Vepefos
35805433|T121|Vepeside
35805434|T121|Vepsid
35805435|T121|Vepside
35805436|T121|Advacan
35805437|T121|Afinitor
35805438|T121|Afinitor Disperz
35805439|T121|Certican
35805378|T121|Everecan
35805379|T121|EverGraf
35805440|T121|Evermil
35805441|T121|Evertor
35805442|T121|Rapact
35805443|T121|Rolimus
35805444|T121|Votubia
35805445|T121|Zortress
35805446|T121|EVAIA
35805446|T121|Etoposide, Vincristine, Adriamycin (Doxorubicin), Ifosfamide, DActinomycin
35805447|T121|VACA
35805447|T121|Vincristine, Adriamycin (Doxorubicin), Cyclophosphamide, DActinomycin
912064|T121|ddAC and Atezolizumab
912064|T121|dose-dense Adriamycin (Doxorubicin), Cyclophosphamide, Atezolizumab
35805448|T121|VACA/IE
35805448|T121|Vincristine, Adriamycin (Doxorubicin), Cyclophosphamide, DActinomycin alternating with Ifosfamide, Etoposide
35805449|T121|VAIA
35805449|T121|Vincristine, Adriamycin (Doxorubicin), Ifosfamide, Actinomycin-D (Dactinomycin)
35805450|T121|VDC/IE
35805450|T121|VAdriaC/IE
35805450|T121|Vincristine, Doxorubicin, Cyclophosphamide, alternating with Ifosfamide and Etoposide
35805450|T121|Vincristine, Adriamycin (Doxorubicin), Cyclophosphamide, alternating with Ifosfamide and Etoposide
912065|T121|Targeted therapy
35805451|T121|VIDE
35805451|T121|Vincristine, Ifosfamide, Doxorubicin, Etoposide
35805452|T121|VAI
35805452|T121|IVA
35805452|T121|Vincristine, DActinomycin, Ifosfamide
35805452|T121|Ifosfamide, Vincristine, DActinomycin
35805452|T121|Vincristine, Actinomycin-D (Dactinomycin), Ifosfamide
35805452|T121|Ifosfamide, Vincristine, Actinomycin-D (Dactinomycin)
35805453|T121|Cyclophosphamide and Topotecan
912066|T121|TG plus Bev
35805454|T121|IE
35805454|T121|Ifosfamide, Etoposide
35805454|T121|Ifosfamide and Etoposide
912067|T121|TH (Taxol) and Everolimus
35805455|T121|Irinotecan and Temozolomide
35805456|T121|TC, then IE, VDoxoC, VEC
35805456|T121|Topotecan, Cyclophosphamide followed by Ifosfamide, Etoposide, then Vincristine, Doxorubicin, Cyclophosphamide, then Vincristine, Etoposide, Cyclophosphamide
35805457|T121|VAdCA
35805457|T121|Vincristine, Adriamycin (Doxorubicin), Cyclophosphamide, DActinomycin
35805458|T121|VAdCA/IE
35805458|T121|Vincristine, Adriamycin (Doxorubicin), Cyclophosphamide, DActinomycin alternating with Ifosfamide, Etoposide
35805459|T121|Aromadex
35805460|T121|Aromasin
35805461|T121|Aromex
35805462|T121|Xtane
35805463|T121|DEP and RT
35805463|T121|Dexamethasone, Etoposide, Platinol (Cisplatin), Radiation Therapy
35805464|T121|DeVIC and RT
35805464|T121|Dexamethasone, VP-16 (Etoposide), Ifosfamide, Carboplatin, Radiation Therapy
912068|T121|TMB-H
35805465|T121|GELOX/RT
35805465|T121|Gemcitabine, L-asparaginase, Oxaliplatin, alternating with Radiation Therapy
35805466|T121|LVP .22Sandwich.22
35805466|T121|LVP
35805466|T121|L-asparaginase, Vincristine, Prednisolone
35805467|T121|MESA/RT
35805467|T121|Methotrexate, Etoposide, Steroid (dexamethasone), PEG-A-sparaginase alternating with Radiation Ttherapy
912069|T121|TP
35805468|T121|SMILE
35805468|T121|Steroid (Dexamethasone), Methotrexate, Ifosfamide, L-asparaginase, Etoposide
35805469|T121|AspaMetDex
35805469|T121|Asparaginase, Methotrexate, Dexamethasone
912070|T121|Trifluridine and tipiracil and Bevacizumab
912071|T121|trimetrexate glucuronate
912071|T121|Trimetrexate
35805470|T121|Alphanine SD
35805471|T121|Mononine
35805472|T121|BeneFix
35805473|T121|Alprolix
35805474|T121|Hemofil-M
35805475|T121|Koate-DVI
35805476|T121|Koate-HP
35805477|T121|Monarc-M
35805478|T121|Monoclate-P
35805479|T121|Advate rAHF-PFM
35805480|T121|Helixate
35805481|T121|Helixate FS
35805482|T121|Kogenate
35805483|T121|Kogenate FS
35805484|T121|Recombinate
35805485|T121|Refacto
35805486|T121|Xyntha
35805487|T121|AryoSeven
35805488|T121|NovoSeven
35805489|T121|NovoSeven RT
35805490|T121|Novo-Seven
35805491|T121|NovoSeven room temperature stable
35805492|T121|Factor X human
35805493|T121|Coagadex
35805494|T121|Corifact
35805495|T121|Famvir
35805496|T121|Pepcid
35805497|T121|Injectafer
35805498|T121|Ferrlecit
35805499|T121|Fe Tabs
35805500|T121|Feosol
35805501|T121|Fer Iron
35805502|T121|Fer-Gen-Sol
35805503|T121|Fer-in-Sol
35805504|T121|Fer-Iron
35805505|T121|Feratab
35805506|T121|FeroSul
35805507|T121|Ferra-TD
35805508|T121|Ferra T.D. Caps
35805509|T121|Ferro-Bob
35805510|T121|Feraheme
35805511|T121|Zarxio
35805512|T121|Biocilin
35805513|T121|Biofigran
35805514|T121|Biofilgran
35805515|T121|Euprotin
35805516|T121|Filatil
35805517|T121|Filgen
35805518|T121|Filgrastima
35805519|T121|Gran
35805520|T121|Granulokine
35805521|T121|Grasalva
35805522|T121|Grasin
35805523|T121|Grastim
35805524|T121|Leicita
35805525|T121|Leubene
35805526|T121|Leucin
35805527|T121|Leucocim
35805528|T121|Leucokain
35805529|T121|Leucostim
35805530|T121|Leukokine
35805531|T121|Leumostin
35805532|T121|Lioplim
35805533|T121|Mielastra
35805534|T121|Myelostim
35805535|T121|Neipogen
35805536|T121|Neitrostim
35805537|T121|Neukine
35805538|T121|Neupogen
35805539|T121|Nevkine
35805540|T121|Nivestim
35805541|T121|Topneuter
35805542|T121|Proscar
35805543|T121|FUDF
35805544|T121|Diflucan
35805545|T121|Beneflur
35805546|T121|Fludabine
35805547|T121|Fludara
35805548|T121|Lymfuda
35805549|T121|Oforta
35805550|T121|Accusite
35805551|T121|Actino Hermal
35805552|T121|Adrucil
35805553|T121|Arumel
35805554|T121|Benton
35805555|T121|Biofur
35805556|T121|Carac
35805557|T121|Carebin
35805558|T121|Carzonal
35805559|T121|Cinco-FU
35805560|T121|Cinkef-U
35805561|T121|Curacil
35805562|T121|Effcil
35805563|T121|Efudex
35805564|T121|Efurix
35805565|T121|Ezadex
35805566|T121|Fauldfluor
35805567|T121|Fivocil
35805568|T121|Fivoflu
35805569|T121|Flacule
35805570|T121|Flonida
35805571|T121|Florac
35805572|T121|Fluhomer
35805573|T121|Fluolex
35805574|T121|Fluoroplex
35805575|T121|Fluor-Uracil
35805576|T121|Fluoro-Uracile ICN
35805577|T121|Fluoro-Uracil ICN
35805578|T121|Fluorouracile
35805579|T121|Fluorouracilo
35805580|T121|Fluorourcil
35805581|T121|Fluoruracilo
35805582|T121|Fluoxan
35805583|T121|Flurablastin
35805584|T121|Flurac
35805585|T121|Fluracedyl
35805586|T121|Fluracil
35805587|T121|Fluroblastin
35805588|T121|Fluroblastine
35805589|T121|Ftoruracil
35805590|T121|Ftouracil
35805591|T121|Haemato-FU
35805592|T121|Ifacil
35805593|T121|Kang Ning
35805594|T121|Kecimeton Tatumi
35805595|T121|Killit
35805596|T121|Lunachol
35805597|T121|Lunapon
35805598|T121|Natira U
35805599|T121|Neofluor
35805600|T121|O Fluor
35805601|T121|Oncofu
35805602|T121|Onkofluor
35805603|T121|Pentafu
35805604|T121|Pharmauracil
35805605|T121|Phthoruracil
35805606|T121|Phtoruracil
35805607|T121|Ribofluor
35805608|T121|Rotianin
35805609|T121|Satelol
35805610|T121|Seco Uracil
35805611|T121|Tecflu
35805612|T121|Timadin
35805613|T121|Triosules
35805614|T121|Uflahex
35805615|T121|Ulosagen
35805616|T121|Ulup
35805617|T121|Uraciflor
35805618|T121|Utoral
35805619|T121|Vaflu
35805620|T121|Vafu
35805621|T121|Halotestin
35805622|T121|Ultandren
35805623|T121|Cytomid
35805624|T121|Eulexin
35805625|T121|Flutamid
35805626|T121|Flutatec
35805627|T121|Lutamide
35805628|T121|Proscan
35805629|T121|Tamid
912072|T121|TX plus Bev
35805630|T121|R-CVP
35805630|T121|Rituximab, Cyclophosphamide, Vincristine, Prednisone
35805631|T121|Rituximab monotherapy, extended course
35805632|T121|Rituximab monotherapy, very extended course
912073|T121|Vinorelbine and Trastuzumab (VH) and Everolimus
912073|T121|VH and Everolimus
912073|T121|Vinorelbine, Herceptin (Trastuzumab), Everolimus
35805633|T121|G-CVP
35805633|T121|Gazyva (Obinutuzumab), Cyclophosphamide, Vincristine, Prednisone
35805634|T121|G-CHOP
35805634|T121|Gazyva (Obinutuzumab), Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
35805635|T121|Rituximab monotherapy, abbreviated course
912074|T121|TX-CEX
912074|T121|Taxotere (Docetaxel) and Xeloda (Capecitabine) followed by Cyclophosphamide, Epirubicin, Xeloda (Capecitabine)
35805636|T121|R-CHVP plus I
35805636|T121|R-CHVP+I
35805636|T121|Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), VP-16 (Etoposide), Prednisolone, Interferon-a2a
35805637|T121|Interferon alfa-2a monotherapy
35805638|T121|R-FM
35805638|T121|FMR
35805638|T121|Rituximab, Fludarabine, Mitoxantrone
35805638|T121|Fludarabine, Mitoxantrone, Rituximab
35805639|T121|R-FND
35805639|T121|Rituximab, Fludarabine, Novantrone (mitoxantrone), Dexamethasone
35805639|T121|Rituximab, Fludarabine, Novantrone, Dexamethasone
35805640|T121|O-CHOP
35805640|T121|Ofatumumab, Cyclophosphamide, Hydroxydaunorubicin, Oncovin, Prednisone
35805641|T121|R-CMD
35805641|T121|Rituximab, Cladribine, Mitoxantrone, Dexamethasone
35805642|T121|Bortezomib and Rituximab (VR)
35805642|T121|VR
35805642|T121|Velcade (Bortezomib) and Rituximab
35805642|T121|Velcade (Bortezomib), Rituximab
35805643|T121|FM
35805643|T121|Fludarabine, Mitoxantrone
35805645|T121|Bevacizumab and Rituximab
35805646|T121|BVR
35805646|T121|VBR
35805646|T121|Bendamustine, Velcade (Bortezomib), Rituximab
35805646|T121|Velcade (Bortezomib), Bendamustine, Rituximab
35805647|T121|Copanlisib monotherapy
35805648|T121|Lenalidomide, Dexamethasone, Rituximab
35805649|T121|PEP-C
35805649|T121|Prednisone, Etoposide, Procarbazine, Cyclophosphamide
35805650|T121|Vorinostat and Rituximab
35805651|T121|VR-CP
35805651|T121|Velcade (Bortezomib), Rituximab, Cyclophosphamide, Prednisone
35805652|T121|FCR, then allo HSCT
35805652|T121|Fludarabine, Cyclophosphamide, Rituximab
35805644|T121|(90)YFC, then allo HSCT
35805644|T121|Ibritumomab tiuxetan, Fludarabine, Cyclophosphamide
35805653|T121|CHOP, then 131Iodine-Tositumomab
35805653|T121|CHOP-RIT
35805653|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne RadioImmunoTherapy
35805654|T121|CHVP
35805654|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Vumon (Teniposide), Prednisone
35805654|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Vm26 (Teniposide), Prednisone
35805655|T121|CHVP-I
35805655|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Vumon (Teniposide), Prednisone, Interferon alfa-2b
35101760|T121|Baklinger
35805656|T121|COPA
35805656|T121|Cyclophosphamide, Oncovin (Vincristine), Prednisone, Adriamycin (Doxorubicin)
912075|T121|MSC-2156119
912075|T121|EMD-1214063
912075|T121|MSC-2156119J
912075|T121|Tepotinib
35101759|T121|Baktar
35101758|T121|Bakton
35101757|T121|Baktrisid DS
35805657|T121|CVP, then 131Iodine-Tositumomab
35805657|T121|CVP-RIT
35805657|T121|Cyclophosphamide, Vincristine, Prednisone, then RadioImmunoTherapy
35805658|T121|Fludarabine, then 131Iodine-Tositumomab
35805659|T121|FND
35805659|T121|Fludarabine, Novantrone (Mitoxantrone), Dexamethasone
35805660|T121|131Iodine-Tositumomab monotherapy
35805661|T121|MCP
35805661|T121|Mitoxantrone, Chlorambucil, Prednisone
35805662|T121|FMP
35805662|T121|Fludarabine, Mitoxantrone, Prednisone
35805663|T121|Arixtra
35805664|T121|Quixidar
35805665|T121|Fodosine
35805666|T121|Mundesine
35805667|T121|Emend for Injection
35805668|T121|Tavalisse
35805669|T121|Muphoran
35805670|T121|Mustophoran
35805671|T121|Faslodex
35805672|T121|Fasnorm
35805673|T121|Fulvenat
35805674|T121|Fulvidax
35805675|T121|Fuvestrol
35805676|T121|Lasix
35805677|T121|Salix
35805678|T121|Gastrectomy
35101756|T121|Balkatrin
35101755|T121|Balkatrine
35805679|T121|FP/Capecitabine and RT
35805679|T121|Fluorouracil and Platinol (Cisplatin) alternating with Capecitabine and Radiation Therapy
912076|T121|Doxorubicin, L-asparaginase, Mercaptopurine, Vincristine, Prednisone
35805680|T121|Cisplatin and S-1
35805680|T121|CS
35805680|T121|SP
35805680|T121|S-1 and Platinol (Cisplatin)
912077|T121|EC-D
912077|T121|Epirubicin and Cyclophosphamide followed by Docetaxel
912077|T121|Epirubicin and Cyclophosphamide followed by Taxotere (Docetaxel)
912078|T121|Epoetin beta
35805681|T121|Docetaxel and S-1
35805681|T121|DS
912079|T121|Flagyl
912080|T121|Fludarabine and TBI for haploidentical transplant
912080|T121|Flu/TBI
912080|T121|<u><b>Flu</b></u>darabine and Total Body Irradiation
35805682|T121|Fluorouracil, Folinic acid, Mitomycin
35805683|T121|OLF
35805683|T121|FLO
35805683|T121|Oxaliplatin, Leucovorin, Fluorouracil
35805683|T121|Fluorouracil, Leucovorin, Oxaliplatin
35805683|T121|OFF
35805683|T121|Oxaliplatin, Leucovorin (Folinic acid), Fluorouracil
35805683|T121|Oxaliplatin, Fluorouracil, Folinic acid
35805684|T121|Paclitaxel and S-1
35805685|T121|UFTM
35805685|T121|UFT (Tegafur and uracil) and Mitomycin
912081|T121|Cisplatin and Gemcitabine (GC) and Atezolizumab
912081|T121|GC and Atezolizumab
912081|T121|Gemcitabine, Cisplatin, Atezolizumab
912082|T121|Carboplatin and Gemcitabine (GCb) and Atezolizumab
912082|T121|GCb and Atezolizumab
912082|T121|Gemcitabine, Carboplatin, Atezolizumab
35805686|T121|Doxifluridine and Mitomycin
35805687|T121|FAM
35805687|T121|Fluorouracil, Adriamycin (Doxorubicin), Mitomycin
35805688|T121|FAMTX
35805688|T121|Fluorouracil, Adriamycin (Doxorubicin), MTX (Methotrexate)
35805689|T121|FEMTX
35805689|T121|Fluorouracil, Epirubicin, MTX (Methotrexate)
35805690|T121|Pazopanib monotherapy
35805691|T121|Sunitinib monotherapy
35805692|T121|Cangib
35805693|T121|Denrit
35805694|T121|Geffy
35805695|T121|Gefitec
35805696|T121|Gefitero
35805697|T121|Gefonib
35805698|T121|Geftib
35805699|T121|Geftican
35805700|T121|Gefticip
35805701|T121|Geftilon
35805702|T121|Geftinat
35805703|T121|Geftiwel
35805704|T121|Iressa
35805705|T121|KabiGef
35805706|T121|Gemcite
35805707|T121|Gemzar
35805708|T121|Mylotarg
35805709|T121|Xospata
35805710|T121|Daurismo
35805711|T121|Bevacizumab and RT
35805711|T121|Bevacizumab and Radiation Therapy
35805712|T121|Carmustine and RT
35805712|T121|BCNU and RT
35805712|T121|BCNU (Carmustine) and Radiation Therapy
35805713|T121|Nimustine and RT
35805713|T121|Nimustine and Radiation Therapy
35101754|T121|Bantizol
35805714|T121|Temozolomide and low-dose RT
35805714|T121|Temozolomide and LDRT
35805714|T121|Temozolomide and Low-Dose Radiation Therapy
35805715|T121|Temozolomide and NovoTTF-100A
35805716|T121|PMA P100034/S013
35805716|T121|NovoTTF-100A system (Optune)
35805717|T121|Gliadel wafer monotherapy
912083|T121|Inqovi
35805718|T121|Hydroxyurea and Imatinib
35805719|T121|Lomustine monotherapy
35805720|T121|NovoTTF-100A monotherapy
35805721|T121|Voraxaze
35805722|T121|Novgos
35805723|T121|Zoladex
35805724|T121|Prophylaxis
35805725|T121|Cyclosporine and Methotrexate
35805726|T121|Cyclosporine, Methotrexate, ATG
35805727|T121|Cyclosporine, Methotrexate, Methylprednisolone
35805728|T121|Cyclosporine, Methotrexate, Prednisone
35805729|T121|Methotrexate, Tacrolimus, Tocilizumab
35805730|T121|Methotrexate, Tacrolimus, Vorinostat
35805731|T121|Rabbit ATG
35805732|T121|Cyclosporine and Prednisone
35805733|T121|Cyclosporine, Corticosteroids, Rituximab
35805734|T121|Cyclosporine, Sirolimus, Prednisone
35805735|T121|Sirolimus, Tacrolimus, Prednisone
35805736|T121|Gramatic
35805737|T121|Granicip
35805738|T121|Graniset
35805739|T121|Granisev
35805740|T121|Granisol
35805741|T121|Granitero
35805742|T121|Graniz
35805743|T121|Granney
35805744|T121|Granny
35805745|T121|Granovell
35805746|T121|Gratryl
35805747|T121|Kytril
35805748|T121|Naurif
35805749|T121|Sancuso
35805750|T121|Sustol
35805751|T121|dmCODOX-M - Modified Magrath
35805751|T121|dmCODOX-M
35805751|T121|dose-modified Cyclophosphamide, Oncovin, DOXorubicin, Methotrexate
35805752|T121|dmCODOX-M/IVAC - Modified Magrath
35805752|T121|dmCODOX-M/IVAC
35805752|T121|dose-modified Cyclophosphamide, Oncovin, DOXorubicin, Methotrexate alternating with Ifosfamide, Vepesid (etoposide), Ara-C (cytarabine)
35805753|T121|EPOCH, dose-escalated
35805753|T121|Etoposide, Prednisone, Oncovin (Vincristine), Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin)
35805754|T121|R-EPOCH, dose-escalated
35805754|T121|Rituximab, Etoposide, Prednisone, Oncovin (Vincristine), Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin)
35805755|T121|SC-EPOCH-RR
35805755|T121|Short Course Rituximab, Etoposide, Prednisone, Oncovin, Cyclophosphamide, Hydroxydaunorubicin, with dose-dense Rituximab
35805756|T121|Stanford V
912084|T121|Liso-cel
912085|T121|JCAR017
912085|T121|Lisocabtagene maraleucel
35805757|T121|Cladribine and Rituximab
912086|T121|MAC
912086|T121|Mitoxantrone and Ara-C (Cytarabine)
912086|T121|Mitoxantrone and Intermediate-Dose Ara-C (Cytarabine)
35805758|T121|Moxetumomab pasudotox monotherapy
35805759|T121|Haldol
35805760|T121|Heloper
35805761|T121|Serenace
35805762|T121|Trancodol
35805763|T121|Laryngectomy
35805764|T121|Head and neck cancer surgery
35805765|T121|No induction
35805766|T121|Cetuximab and RT
35805766|T121|Cetuximab and Radiation Therapy
35805767|T121|Carboplatin, Fluorouracil, Cetuximab, RT
35805767|T121|Carboplatin, Fluorouracil, Cetuximab, Radiation Therapy
35805768|T121|Docetaxel, Fluorouracil, Hydroxyurea, RT
35805768|T121|DFHX
35805768|T121|Docetaxel, Fluorouracil, Hydroxyurea, XRT (Radiation therapy)
35805769|T121|Fluorouracil, Hydroxyurea, RT
35805769|T121|Fluorouracil, Hydroxyurea, Radiation Therapy
35805770|T121|Cisplatin, Cetuximab, RT
35805770|T121|Cisplatin, Cetuximab, Radiation Therapy
35805771|T121|Docetaxel, Cetuximab, RT
35805771|T121|Docetaxel, Cetuximab, Radiation Therapy
35805772|T121|Tegafur and Uracil
35805773|T121|Carboplatin and Fluorouracil
35805774|T121|Carboplatin, Fluorouracil, Cetuximab
35805775|T121|Cisplatin and Cetuximab
35805776|T121|Cisplatin and Fluorouracil (CF) and Panitumumab
35805777|T121|Bleomycin, Methotrexate, Vinblastine/RT
35805778|T121|CABO
35805778|T121|Cisplatin, Amithopterin (Methotrexate), Bleomycin, Oncovin (Vincristine)
35805779|T121|Hemacord
35805780|T121|HLH-94 regimen
35805781|T121|Antifungals
35805782|T121|HLH-2004 regimen
35805783|T121|IVIG
35805783|T121|Intravenous immunoglobulin
35805784|T121|DEP
35805784|T121|Doxil (Pegylated liposomal doxorubicin), Etoposide, MethylPrednisolone
35805785|T121|Argatroban monotherapy
35805786|T121|Danaparoid monotherapy
35805787|T121|Fondaparinux monotherapy
35805788|T121|Lepirudin monotherapy
35805789|T121|Axitinib and TACE
35805790|T121|TACE
35805791|T121|DEB-TACE
35805791|T121|Drug-Eluting Bead Trans-Arterial Chemo-Embolization
35805792|T121|Radioembolization
35805793|T121|TACE monotherapy
35805793|T121|Trans-Arterial Chemo-Embolization
35805794|T121|Hepatobiliary cancer surgery
35101753|T121|Basatin
35805795|T121|Lenvatinib monotherapy
35805796|T121|TACE, then 5-FU
35805796|T121|Trans-Arterial ChemoEmbolization followed by 5-FluoroUracil
35101752|T121|Baserin
35805797|T121|Cabozantinib monotherapy
35805798|T121|SunPla
35805799|T121|Tamoxifen acid monotherapy
35805800|T121|Tranexamic acid monotherapy
35805801|T121|Vantas
35805802|T121|ABVD
35805802|T121|Adriamycin (Doxorubicin), Bleomycin, Vinblastine, Dacarbazine
35805803|T121|eBEACOPP
35805803|T121|escalated Bleomycin, Etoposide, Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Procarbazine, Prednisone
35805803|T121|escBEACOPP
35805803|T121|BEACOPP(escalated)
35805803|T121|Bleomycin, Etoposide, Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Procarbazine, Prednisone, escalated dose
35805804|T121|AVD
35805804|T121|Adriamycin (Doxorubicin), Vinblastine, Dacarbazine
35805805|T121|MOPP-ABV
35805805|T121|Mustargen (Mechlorethamine), Oncovin (Vincristine), Procarbazine, Prednisone, Adriamycin (Doxorubicin), Bleomycin, Vinblastine
35805806|T121|VAMP (Methotrexate)
35805806|T121|Vinblastine, Adriamycin (Doxorubicin), Methrotrexate, Prednisone
35805807|T121|A-AVD
35805807|T121|A+AVD
35805807|T121|BV + AVD
35805807|T121|Adcetris (Brentuximab vedotin), Adriamycin (Doxorubicin), Vinblastine, Dacarbazine
35805807|T121|Brentuximab Vedotin, Adriamycin (Doxorubicin), Vinblastine, Dacarbazine
35805807|T121|B-AVD
35805807|T121|AVD-A
35805807|T121|Brentuximab vedotin, Adriamycin (Doxorubicin), Vinblastine, Dacarbazine
35805807|T121|Adriamycin (Doxorubicin), Vinblastine, Dacarbazine, Adcetris (Brentuximab vedotin)
35805808|T121|BEACOPP
35805808|T121|Bleomycin, Etoposide, Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Procarbazine, Prednisone
35805808|T121|bBEACOPP
35805808|T121|baseline Bleomycin, Etoposide, Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Procarbazine, Prednisone
35805809|T121|EBVP
35805809|T121|Epirubicin, Bleomycin, Vinblastine, Prednisone
35805810|T121|RABVD
35805810|T121|Rituximab, Adriamycin (Doxorubicin), Bleomycin, Vinblastine, Dacarbazine
35805811|T121|IGEV
35805811|T121|Ifosfamide, GEmcitabine, Vinorelbine
35805812|T121|BEACOPP-14
35805812|T121|Bleomycin, Etoposide, Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine), Procarbazine, Prednisone, 14-day course
35805813|T121|ABVD, DD-DI
35805813|T121|Adriamycin (Doxorubicin), Bleomycin, Vinblastine, Dacarbazine, Dose-Dense and Dose-Intense
912087|T121|Hematologic monoclonal antibody
35805814|T121|C-MOPP/ABV
35805814|T121|CyclophosphaMide, Oncovin (Vincristine), Procarbazine, Prednisone, Adriamycin (Doxorubicin), Bleomycin, Vinblastine
35805815|T121|MOPP
35805815|T121|Mechlorethamine, Oncovin (Vincristine), Procarbazine, Prednisone
35101751|T121|Batrox
35805816|T121|VEBEP
35805816|T121|Vepesid (Etoposide), Epirubicin, Bleomycin, Endoxan (Cyclophosphamide), Prednisolone
35805817|T121|ABVE-PC
35805817|T121|Adriamycin (Doxorubicin), Bleomycin, Vincristine, Etoposide, Prednisone, Cyclophosphamide
35805818|T121|OEPA
35805819|T121|COPDAC
35805819|T121|Cyclophosphamide, Oncovin (Vincristine), Prednisone, DACarbazine
35805820|T121|OPPA
35805820|T121|Oncovin (Vincristine), Procarbazine, Prednisone, Adriamycin (Doxorubicin)
35805821|T121|Brentuximab vedotin and Dacarbazine
35805822|T121|ChlVPP
35805822|T121|Chllorambucil, Vinblastine, Procarbazine, Prednisone
35805823|T121|ChlVPP/EVA
35805823|T121|Chllorambucil, Vinblastine, Procarbazine, Prednisone, Etoposide, Vincristine, Adriamycin (Doxorubicin)
35805824|T121|PVAG
35805824|T121|Prednisone, Vinblastine, Adriamycin (Doxorubicin), Gemcitabine
35805825|T121|VEPEMB
35805825|T121|Vinblastine, Endoxan (Cyclophosphamide), Procarbazine, Etoposide, Mitoxantrone, Bleomycin
35805826|T121|COPP/ABVD
35805826|T121|C-MOPP/ABVD
35805826|T121|Cyclophosphamide, Oncovin (Vincristine), Procarbazine, Prednisone alternating with Adriamycin (Doxorubicin), Bleomycin, Vinblastine, Dacarbazine
35805826|T121|CyclophosphaMide, Oncovin (Vincristine), Procarbazine, Prednisone alternating with Adriamycin (Doxorubicin), Bleomycin, Vinblastine, Dacarbazine
35805827|T121|BeGEV
35805827|T121|Bendamustine, GEmcitabine, Vinorelbine
35805828|T121|Brentuximab vedotin and Nivolumab
35805829|T121|BVB
35805830|T121|DexaBEAM
35805830|T121|Dexamethasone, BiCNU (Carmustine), Etoposide, Ara-C (Cytarabine), Melphalan
35805831|T121|DHAP - time intensified
35805831|T121|Dexamethasone, High-dose Ara-C (Cytarabine), Platinol (Cisplatin)
35805832|T121|GCD
35805832|T121|Gemcitabine, Carboplatin, Dexamethasone
35805833|T121|GCD-R
35805833|T121|Gemcitabine, Carboplatin, Dexamethasone, Rituximab
35805834|T121|Gemcitabine and Rituximab
35805834|T121|R-G
35805834|T121|Rituximab and Gemcitabine
35805835|T121|GVP
35805835|T121|Gemcitabine, Vinorelbine, Prednisolone
35805836|T121|Ifosfamide and Vinorelbine
35805837|T121|Mini-BEAM
35805837|T121|dose-reduced BiCNU (Carmustine), Etoposide, Ara-C (Cytarabine), Melphalan
35805838|T121|O-ESHAP
35805838|T121|Ofatumumab, Etoposide, Solumedrol (Methylprednisolone) High-dose Ara-C (Cytarabine), Platinol (Cisplatin)
35101750|T121|Baxolex
35805839|T121|Vinblastine monotherapy
35805840|T121|CBV-Mx, then auto HSCT
35805841|T121|Flu-Mel, then allo HSCT
35805841|T121|Flu-Mel
35805842|T121|Fludarabine, Melphalan, Alemtuzumab, then allo HSCT
35805843|T121|ABVDm
35805843|T121|Adriamycin (Doxorubicin), Bleomycin, Vinblastine, Dacarbazine, methylprednisolone
35805844|T121|BCVPP
35805844|T121|BCNU (Carmustine), Cyclophosphamide, Vincristine, Procarbazine, Prednisone
35805845|T121|ChlVPP/PABIOE
35805845|T121|Chlorambucil, Vinblastine, Procarbazine, Prednisone alternating with Prednisolone, Adriamycin (Doxorubicin), Bleomycin, Oncovin (Vincristine), Etoposide
35101749|T121|bb2121
35101749|T121|ide-cel
35101749|T121|Idecabtagene vicleucel
35805846|T121|COPP (CCNU)
35805846|T121|COPP
35805846|T121|CCNU (Lomustine), Oncovin (Vincristine), Procarbazine, Prednisone
35805847|T121|CVPP
35805847|T121|CCNU (Lomustine), Vinblastine, Procarbazine, Prednisone
35805848|T121|Doxorubicin and Vinblastine
35805849|T121|LOPP
35805849|T121|Leukeran (Chlorambucil), Oncovin (Vincristine), Procarbazine, Prednisone
35805850|T121|LOPP/EVAP
35805850|T121|Leukeran (Chlorambucil), Oncovin (Vincristine), Procarbazine, Prednisone alternating with Etoposide, Vinblastine, Adriamycin (Doxorubicin), Prednisone
35805851|T121|Mechlorethamine monotherapy
35805852|T121|MOPP/ABVD
35805852|T121|Mustargen (Mechlorethamine), Oncovin (Vincristine), Procarbazine, Prednisone alternating with Adriamycin (Doxorubicin), Bleomycin, Vinblastine, Dacarbazine
35805853|T121|MVPP
35805853|T121|Mechlorethamine, Vinblastine, Procarbazine, Prednisone
35805854|T121|NOVP
35805854|T121|Novantrone (Mitoxantrone), Oncovin (Vincristine), Vinblastine, Prednisone
35805855|T121|SCAB
35805855|T121|Streptozocin, CCNU (Lomustine), Adriamycin (Doxorubicin), Bleomycin
35805856|T121|ABDIC
35805856|T121|Adriamycin (Doxorubicin), Bleomycin, DIC (Dacarbazine), CCNU (Lomustine), Prednisone
35805857|T121|B-CAVe
35805857|T121|Bleomycin, CCNU (Lomustine), Adriamycin (Doxorubicin), Vinblastine
35805858|T121|BVCPP
35805858|T121|BCNU (Carmustine), Vinblastine, Cyclophosphamide, Procarbazine, Prednisone
35805859|T121|BVDS
35805859|T121|Bleomycin, Vinblastine, Doxorubicin, Streptozocin
35805860|T121|CEP
35805860|T121|CCNU (Lomustine), Etoposide, Prednimustine
35805860|T121|Cyclophosphamide, Epirubicin, Platinol (Cisplatin)
35805861|T121|CVB
35805861|T121|CCNU (Lomustine), Vinblastine, Bleomycin
35805862|T121|Doxorubicin and Lomustine
35805863|T121|Sirolimus and Vorinostat
35805864|T121|Cortef
35805865|T121|Biosupressin
35805866|T121|Cytodrox
35805867|T121|Droxia
35805868|T121|Droxiurea
35805869|T121|Durea
35805870|T121|Hidrea
35805871|T121|Hondrea
35805872|T121|Hydab
35805873|T121|Hydrea
35805874|T121|Hydrine
35805875|T121|Hydrourea
35805876|T121|Hytas
35805877|T121|Litalir
35805878|T121|Myelostat
35805879|T121|Mylocel
35805880|T121|Neodrea
35805881|T121|Onco Carbide
35805882|T121|Siklos
35805883|T121|Syrea
35805884|T121|Ureax
35805885|T121|Cladribine and Cytarabine
35805886|T121|Mepolizumab monotherapy
35805887|T121|Bandrobon
35805888|T121|Bandrone
35805889|T121|Bondenza
35805890|T121|Bondronat
35805891|T121|Bonviva
35805892|T121|Femorel
35805893|T121|Zevalin
35805894|T121|Imbruvica
35805895|T121|Conmana
35805896|T121|Idamycin
35805897|T121|Idaru
35805898|T121|Ondarubin
35805899|T121|Zavedos
35805900|T121|Zavedose
35805901|T121|Praxbind
35805902|T121|Zydelig
35805903|T121|Enliven
35805904|T121|Glivec
35805905|T121|Gleevac
35805906|T121|Gleevec
35805907|T121|Imalek
35805908|T121|Imatib
35805909|T121|Temsan
35805910|T121|Veenat
35805911|T121|Dexamethasone and Eltrombopag
35805913|T121|Dexamethasone and Rituximab
35805914|T121|Intravenous immunoglobulin monotherapy
35805914|T121|IntraVenous ImmunoGlobulin
35805915|T121|RhIG monotherapy
35805915|T121|RhIG
35805915|T121|Rho(D) Immune Globulin
35805916|T121|TT4
35805916|T121|Triple Therapy (4?)
35805917|T121|ATRA and Danazol
35805918|T121|Avatrombopag monotherapy
35805919|T121|Danazol monotherapy
35805920|T121|Fostamatinib monotherapy
35805921|T121|Mycophenolate mofetil monotherapy
35805922|T121|Romiplostim monotherapy
35805923|T121|Emicizumab monotherapy
35805924|T121|Besponsa
35805925|T121|Roferon-A
35805926|T121|Flebogamma
35805927|T121|Gammagard
35805928|T121|Gamunex
35805929|T121|Octagam
35805930|T121|Privigen
35805931|T121|Yervoy
35805932|T121|Axinotecan
35805933|T121|Biotecan
35805934|T121|Biskam
35805935|T121|Campto
35805936|T121|Campostar
35805937|T121|Camptosar
35805938|T121|Elinatecan
35805939|T121|Faultenocan
35805940|T121|Irenax
35805941|T121|Irinogen
35805942|T121|Irinotel
35805943|T121|Irinotesin
35805944|T121|Irnocam
35805945|T121|Itoxaril
35805946|T121|Linatecan
35805947|T121|Onivyde
35805948|T121|Satigene
35805949|T121|Tecnotecan
35805950|T121|Tekamen
35805951|T121|Toptecin
35805952|T121|Trinotecan
35805953|T121|Winol
35805954|T121|Dexferrum
35805955|T121|DextraCare
35805956|T121|Ferrodex
35805957|T121|Imferon
35805958|T121|INFeD
35805959|T121|Irondex
35805960|T121|Saferon
35805961|T121|Uniferon
35805962|T121|Venofer
35805963|T121|Accure
35805964|T121|Accutane
35805965|T121|Amnesteem
35805966|T121|Cistane
35805967|T121|Claravis
35805968|T121|Isotrex
35805969|T121|Isotrexin
35805970|T121|Oratane
35805971|T121|Roaccutan
35805972|T121|Roaccutane
35805973|T121|Roacutan
35805974|T121|Sotret
35805975|T121|Sporanox
35805976|T121|Tibsovo
35805977|T121|Ixempra
35805912|T121|Ninlaro
35805978|T121|Nizoral
35805979|T121|Endari
35805980|T121|Epivir
35805981|T121|Etoposide and Prednisone
35805982|T121|Etoposide, Vinblastine, Prednisone
35805983|T121|Methotrexate, Vinblastine, Prednisone
35805984|T121|Vinblastine and Prednisone
35805985|T121|Mercaptopurine, Methotrexate, Vinblastine, Prednisolone
35805986|T121|Ipstyl
35805987|T121|Lanreotide Autogel
35805988|T121|Somatuline Autogel
35805989|T121|Somatuline Depot
35805990|T121|Somatuline LA
35805991|T121|Somatuline LP
35805992|T121|Somatuline PR
35805993|T121|Prevacid
35805994|T121|Tykerb
35805995|T121|Methotrexate and Prednisone
35805996|T121|Vitrakvi
35805997|T121|Kabillon
35805998|T121|Lenalid
35805999|T121|Lenangio
35806000|T121|Lenmid
35806001|T121|Lenome
35806002|T121|Lenzest
35806003|T121|MyeloSar
35806004|T121|Revlimid
35806005|T121|Granocyte
35806006|T121|Neutrogin
35806007|T121|Lenvima
35806008|T121|Refludan
35806009|T121|Femara
35806010|T121|Fempro
35806011|T121|Gynotril
35806012|T121|Latrotal
35806013|T121|Lerozol
35806014|T121|Letoval
35806015|T121|Letpro
35806016|T121|Letromina
35806017|T121|Letroplex
35806018|T121|Letroz
35806019|T121|Letrozol
35806020|T121|Lexel
35806021|T121|Lezole
35806022|T121|Carcinil
35806023|T121|Depo-Eligard
35806024|T121|Eligard
35806025|T121|Enanton
35806026|T121|Enantone
35806027|T121|Enantone-Gyn
35806028|T121|Ginecrin
35806029|T121|Leuplin
35806030|T121|Leupromer
35802850|T121|Leuprorelin
35806031|T121|Leuren
35806032|T121|Lorelin Depot
35806033|T121|Lucrin
35806034|T121|Lucrin Depot
35806035|T121|Lupard Depot
35806036|T121|Lupoide Depot
35806037|T121|Lupride Depot
35806038|T121|Luprodex Depot
35806039|T121|Lupron
35806040|T121|Lupron Depot
35806041|T121|Procren
35806042|T121|Procrin
35806043|T121|Prostap
35806044|T121|Trenantone
35806045|T121|Uno-Enantone
35806046|T121|Valeuprox
35806047|T121|Viadur
35806048|T121|Ergamisol
35806049|T121|Levaquin
35806050|T121|Fusilev
35101748|T121|Befarin
35806051|T121|CRd
35806051|T121|LDC
35806051|T121|RdC
35806051|T121|Cyclophosphamide, Revlimid (Lenalidomide), low-dose dexamethasone
35806051|T121|Lenalidomide, Dexamethasone, Cyclophosphamide
35806051|T121|Revlimid (Lenalidomide), low-dose dexamethasone, Cyclophosphamide
35806051|T121|CLD
35806051|T121|Cyclophosphamide, Lenalidomide Dexamethasone
35806051|T121|Rdc
35806051|T121|Revlimid (Lenalidomide), low-dose dexamethasone, low-dose cyclophosphamide
35806052|T121|Proton pump inhibitors
35806053|T121|Lenalidomide and Dexamethasone (Rd)
35806053|T121|Rd
35806053|T121|RevDex
35806053|T121|Ld
35806053|T121|LenDex
35806053|T121|Revlimid (Lenalidomide) and low-dose dexamethasone
35806053|T121|Revlimid (Lenalidomide) and Dexamethasone
35806053|T121|Lenalidomide and low-dose dexamethasone
35806053|T121|Lenalidomide and Dexamethasone
35806054|T121|CTD
35806054|T121|Cyclophosphamide, Thalidomide, Dexamethasone
35806054|T121|CTDa
35806054|T121|Tdc
35806054|T121|Cyclophosphamide, Thalidomide, Dexamethasone, attenuated
35806054|T121|Thalidomide, low-dose dexamethasone, low-dose cyclophosphamide
35806055|T121|M-DEX
35806055|T121|MD
35806055|T121|Melphalan and DEXamethasone
35806056|T121|Melphalan and Prednisone (MP)
35806056|T121|MP
35806056|T121|Melphalan and Prednisone
35806056|T121|<i>Note
35806056|T121|This regimen is of historical significance</i>
35806057|T121|MRD
35806057|T121|L-M-Dex
35806057|T121|Melphalan, Revlimid (Lenalidomide), Dexamethasone
35806057|T121|Lenalidomide, Melphalan, Dexamethasone
35806058|T121|Melphalan, then auto HSCT
35806059|T121|Bortezomib and Dexamethasone (VD)
35806059|T121|VD
35806059|T121|Velcade (Bortezomib) and D</u>examethasone</b>
35806059|T121|BD
35806059|T121|Velcade (Bortezomib) and Dexamethasone
35806059|T121|Bortezomib and Dexamethasone
35806059|T121|Bd
35806059|T121|Bort-Dex
35806059|T121|Vd
35806059|T121|Velcade (Bortezomib), Dexamethasone
35806059|T121|Bortezomib, Dexamethasone
35806059|T121|Bortezomib, low-dose dexamethasone
35806059|T121|Velcade (Bortezomib), low-dose dexamethasone
35806060|T121|Bortezomib and Melphalan, then auto HSCT
35806061|T121|VDC
35806061|T121|CyBorD
35806061|T121|Velcade (Bortezomib), Dexamethasone, Cyclophosphamide
35806061|T121|Cyclophosphamide, Bortezomib, Dexamethasone
35806061|T121|VDC-mod
35806061|T121|VCD
35806061|T121|Velcade (Bortezomib), Dexamethasone, Cyclophosphamide (modified dose)
35806061|T121|Velcade (Bortezomib), Cyclophosphamide, Dexamethasone
35806061|T121|CVD
35806061|T121|Cyclophosphamide, Velcade (Bortezomib), Dexamethasone
35806062|T121|VMD
35806062|T121|BMDex
35806062|T121|Velcade (Bortezomib), Melphalan, Dexamethasone
35806062|T121|Bortezomib, Melphalan, Dexamethasone
42542277|T121|Acute lymphoblastic leukemia
35806063|T121|Daratumumab monotherapy
35806064|T121|Ixazomib monotherapy
35806065|T121|Ixazomib and Dexamethasone
35806066|T121|Pd
35806067|T121|Lenalidomide and Dexamethasone (RD)
35806067|T121|RD
35806067|T121|Revlimid (Lenalidomide) and high-dose Dexamethasone
35806068|T121|CeeNu
35806069|T121|Gleostine
35806070|T121|Imodium
35806071|T121|Ativan
35806072|T121|Lorbrena
35806073|T121|Carboplatin and Vincristine
35806073|T121|CV
35806073|T121|VC
35806073|T121|Vincristine and Carboplatin
35806074|T121|Carboplatin and Teniposide
35806075|T121|Mulpleta
35806076|T121|Lutathera
35806077|T121|R-DHAC
35806077|T121|Rituximab, Dexamethasone, High-dose Ara-C (Cytarabine), Carboplatin
35806078|T121|R-HiDAC
35806078|T121|Rituximab and High Dose Ara-C (Cytarabine)
35806079|T121|DexaBEAM and G-CSF
35806079|T121|Dexamethasone, BiCNU (Carmustine), Etoposide, Ara-C (Cytarabine), Melphalan, Granulocyte Colony Stimulating Factor
35806080|T121|R-CHOP/R-DHAP
35806080|T121|Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne alternating with Rituximab, Dexamethasone, High-dose Ara-C (Cytarabine), Platinol (Cisplatin)
35806081|T121|Erythrocyte growth factors
42542278|T121|Afatinib and Bevacizumab
35101747|T121|Belfactrin
35806082|T121|VR-CAP
35806082|T121|VcR-CAP
35806082|T121|Velcade (Bortezomib), Rituximab, Cyclophosphamide, Adriamycin (Doxorubicin), Prednisone
42542279|T121|Afatinib and Cetuximab
35806083|T121|maxi-R-CHOP/R-HiDAC
35806083|T121|maximum-strength Rituximab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne alternating with Rituximab, High-Dose Ara-C (Cytarabine)
35806084|T121|TAM6, then auto HSCT
35806085|T121|R-M-CHOP
35806085|T121|Rituximab, MTX (Methotrexate), Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin, Prednisone
35806086|T121|EAR and G-CSF
35806086|T121|Etoposide, Ara-C (Cytarabine), Rituximab, Granulocyte Colony Stimulating Factor
35806087|T121|R-MACLO/R-IVAM
35806087|T121|Rituximab, MTX (Methotrexate), Adriamycin (Doxorubicin), Cyclophosphamide, Leucovorin (Folinic acid), Oncovin (Vincristine) alternating with Rituximab, Ifosfamide, VP-16 (Etoposide), Ara-C (Cytarabine), Mesna
35806088|T121|RiPAD plus C
35806088|T121|RiPAD+C
35806088|T121|Rituximab, PS-341 (Bortezomib), Adriamycin (Doxorubicin), Dexamethasone, Chlorambucil
35806089|T121|R-VAD plus C
35806089|T121|R-VAD+C
35806089|T121|Rituximab, Vincristine, Adriamycin (Doxorubicin), Dexamethasone, Chlorambucil
35806090|T121|Melphalan and TBI, then auto HSCT
35806091|T121|VAD plus C
35806091|T121|VAD+C
35806091|T121|Vincristine, Adriamycin (Doxorubicin), Dexamethasone, Chlorambucil
35806092|T121|VcR-CVAD
35806092|T121|Velcade (Bortezomib), Rituximab, Cyclophosphamide, Vincristine, Adriamycin (Doxorubicin), Dexamethasone
35806093|T121|BCHOP
35806093|T121|Bortezomib, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisolone
35101746|T121|Belon
35806094|T121|Arsenic trioxide and Chlorambucil
35806095|T121|BeRT
35806095|T121|Bendamustine, Rituximab, Temsirolimus
35806096|T121|BDR
35806096|T121|BORID
35806096|T121|Bortezomib, Dexamethasone, Rituximab
35806096|T121|BOrtezomib, RItuximab, Dexamethasone
35806097|T121|Ibrutinib and Venetoclax
35806097|T121|VI
35806097|T121|Ventoclax and Ibrutinib
35806098|T121|RT-PEPC
35806098|T121|Rituximab, Thalidomide, Prednisone, Etoposide, Procarbazine, Cyclophosphamide
35806099|T121|Temsirolimus and Rituximab
35806100|T121|Non-curative second-line consolidation therapy
35806101|T121|BFR, then allo HSCT
35806101|T121|Bendamustine, Fludarabine, Rituximab
35806102|T121|Non-curative second-line maintenance therapy
35806103|T121|Doxycycline monotherapy
35806104|T121|Clarithromycin monotherapy
35101745|T121|Bencole
35806105|T121|Ox-P
35806105|T121|Oxaliplatin and Prednisone
35806106|T121|Chlormethine
35806107|T121|Mustargen
35806108|T121|Mustine
35806109|T121|Depo-Provera
35806110|T121|Provera
35806111|T121|Carboplatin, Cyclophosphamide, Etoposide, Methotrexate, Vincristine
35806112|T121|Cisplatin, Lomustine, Vincristine
35806113|T121|Cyclophosphamide and Vincristine/Cisplatin and Etoposide
35806114|T121|Megace
35806115|T121|CVD, IL-2, IFN alfa-2b - sequential biochemotherapy
35806115|T121|CVD, IL-2, IFN alfa-2b
35806115|T121|bioCT
35806115|T121|Cisplatin, Vinblastine, Dacarbazine, high-dose InterLeukin-2, InterFeroN alfa-2b
35806115|T121|bioChemoTherapy
35806116|T121|Melanoma surgery
35806117|T121|Interferon alfa-2b monotherapy
35806117|T121|HDI
35806117|T121|High-Dose Interferon
35806118|T121|Ipilimumab monotherapy
35101744|T121|Benectrin
35806119|T121|Peginterferon alfa-2b monotherapy
35806120|T121|Lymphadenectomy
912088|T121|Non-small cell lung cancer nonsquamous
912089|T121|Non-small cell lung cancer squamous
35806121|T121|Talimogene laherparepvec monotherapy
35806122|T121|ABC
35806122|T121|Abraxane (Paclitaxel nanoparticle albumin-bound), Bevacizumab, Carboplatin
42542280|T121|BLU-285
42542280|T121|Avapritinib
42542281|T121|Avapritinib monotherapy
35806123|T121|Cisplatin and Dacarbazine
35807525|T121|Cisplatin, Dacarbazine, IL-2, IFN alfa-2b  plus /- Carmustine
35806124|T121|Cisplatin, Dacarbazine, Paclitaxel
35806125|T121|CVD (Vinblastine)
35806125|T121|CVD
35806125|T121|Cisplatin, Vinblastine, Dacarbazine
35806126|T121|CVD (Vindesine)
35806126|T121|CVD
35806126|T121|Cisplatin, Vindesine, Dacarbazine
912090|T121|Panretin
912091|T121|Panretyn
912092|T121|Panrexin
35806127|T121|Dacarbazine monotherapy
42542282|T121|Ayvakit
912093|T121|PLX3397
912093|T121|Pexidartinib
912094|T121|BLU-667
912094|T121|Pralsetinib
912095|T121|Resection
35806128|T121|Dacarbazine and Interferon alfa-2a
35806129|T121|Dacarbazine and Ipilimumab
35806130|T121|Fotemustine monotherapy
35806131|T121|High-dose Interleukin-2
35806131|T121|HD IL-2
35806131|T121|High-Dose InterLeukin-2
35806132|T121|Low-dose Interleukin-2
35806132|T121|LD IL-2
35806132|T121|Low-Dose InterLeukin-2
35806133|T121|Ipilimumab, then Nivolumab
35806134|T121|Nivolumab, then Ipilimumab
35806135|T121|Temozolomide and Bevacizumab
35806135|T121|TB
35806136|T121|IL-2 monotherapy
42542283|T121|BRAF-mutated Melanoma
912096|T121|stilbamidine isetionate
912096|T121|Stilbamidine
912097|T121|Stilbamidine and Urethane
35806137|T121|Binimetinib and Encorafenib
35806138|T121|Cobimetinib and Vemurafenib
912098|T121|Tegafur and uracil monotherapy
35806139|T121|Trametinib monotherapy
35806140|T121|Binimetinib monotherapy
42542284|T121|NRAS-mutated Melanoma
35806141|T121|BCG and Dacarbazine
35806141|T121|BCG and DTIC
35806141|T121|Bacillus Calmette-Guerin and Dimethyl Triazeno Imidazole Carboxamide (Dacarbazine)
35806142|T121|BHD
35806142|T121|BCNU (Carmustine), Hydroxyurea, Dacarbazine
912099|T121|Tumor-reductive surgery
35806143|T121|BVD
35806143|T121|BCNU (Carmustine), Vincristine, Dacarbazine
912100|T121|Turalio
35806144|T121|CDB
35806144|T121|Cisplatin, Dacarbazine, BCNU (Carmustine)
35806145|T121|Cisplatin, Dacarbazine, Interferon alfa-2b
35806146|T121|Cisplatin, Dacarbazine, Tamoxifen
35806147|T121|Dacarbazine and Tamoxifen
35806148|T121|Alkeran
35806149|T121|Alkerana
35806150|T121|Levofolan
35806151|T121|Melfalan
35806152|T121|Bosatria
35806153|T121|Nucala
35806154|T121|Purinethol
35806155|T121|Purixan (oral suspension formulation)
912101|T121|VBM (Vinblastine)
35806156|T121|Anti Uron
35806157|T121|Mesa
35806158|T121|Mesnex
35806159|T121|Mesnil
35806160|T121|Mestian
35806161|T121|Mistabron
35806162|T121|Mistabronco
35806163|T121|Mitexan
35806164|T121|Mucolene
35806165|T121|Neper
35806166|T121|Novacarel
35806167|T121|Siruta
35806168|T121|Uromes
35806169|T121|Uromitexan
35806170|T121|Uroprot
35806171|T121|Varimesna
35806172|T121|Carboplatin and Pemetrexed
35806172|T121|CP
35806172|T121|Carbo-Pem
35806173|T121|Cisplatin and Pemetrexed
35806173|T121|Pem-Cis
35806173|T121|Cis-Pem
35806173|T121|Pemetrexed and Cisplatin
35806173|T121|"<div class=""toccolours"" style=""background-color:#eeeeee"">"
35806173|T121|CPx
35806174|T121|Cisplatin and Raltitrexed
35806175|T121|Cisplatin, Pemetrexed, Bevacizumab
35806175|T121|PCB
35806175|T121|Pemetrexed, Cisplatin, Bevacizumab
35806176|T121|Gemcitabine and Vinorelbine
35806176|T121|VG
35806176|T121|GV
35806176|T121|G+V
35806176|T121|Vinorelbine and Gemcitabine
35806177|T121|Abitrexate
35806178|T121|Alltrex
35806179|T121|Antifolan
35806180|T121|Artrait
35806181|T121|Biometrox
35806182|T121|Biotrexate
35806183|T121|Caditrex
35806184|T121|Cytotrexate
35806185|T121|Ebetrexat
35806186|T121|Emthexat
35806187|T121|Emthexate
35806188|T121|Ervemin
35806189|T121|Farmitrexat
35806190|T121|Fauldmetro
35806191|T121|Folex PFS
35806192|T121|Folitrax
35806193|T121|Hextrate
35806194|T121|Ifamet
35806195|T121|Imutrex
35806196|T121|Ledertrexate
35806197|T121|Ledertrexato
35806198|T121|Lumexon
35806199|T121|Matrex
35806200|T121|Maxtrex
35806201|T121|Medsatrexate
35806202|T121|Merex
35806203|T121|Metex
35806204|T121|Methobax
35806205|T121|Methoblastin
35806206|T121|Methorex
35806207|T121|Methotrexaat
35806208|T121|Methotrexat
35806209|T121|Methotrexato
35806210|T121|Methotrexatum
35806211|T121|Meticil
35806212|T121|Metolate
35806213|T121|Metotressato
35806214|T121|Metotrexate
35806215|T121|Metotrexato
35806216|T121|Metotrexol
35806217|T121|Metrex
35806218|T121|Metrexan
35806219|T121|Metrexato
35806220|T121|Metrotex
35806221|T121|Mexate
35806222|T121|Miantrex CS
35806223|T121|Neometho
35806224|T121|Neotrexate
35806225|T121|Novatrex
35806226|T121|Oncotrex
35806227|T121|O Trexat
35806228|T121|Pharmatrexate
35806229|T121|Remtrex
35806230|T121|Reumatrex
35806231|T121|Rextop
35806232|T121|Rheumatrex
35806233|T121|Tecnomet
35806234|T121|Texate
35806235|T121|Texorate
35806236|T121|Tratoben
35806237|T121|Tremetex
35806238|T121|Trexall
35806239|T121|Trexan
35806240|T121|Trexeron
35806241|T121|Trixilem
35806242|T121|Unitrexate
35806243|T121|Zexate
35806244|T121|Reglan
35806245|T121|Rydapt
35806246|T121|Lyomit
35806247|T121|Mitocin
35806248|T121|Mitocyte
35806249|T121|Mitosol
35806250|T121|Mitozytrex
35806251|T121|Mutamycin
35806252|T121|Lysodren
35806253|T121|Nitrol
35806254|T121|Novantron
35806255|T121|Novantrone
35806256|T121|Poteligeo
35806257|T121|Lumoxiti
35806258|T121|VMP
35806258|T121|Velcade (Bortezomib), Melphalan, Prednisone
35806258|T121|Melphalan, Prednisone, Velcade (Bortezomib)
35806259|T121|VTD
35806259|T121|Velcade (Bortezomib), Thalidomide, Dexamethasone
35806259|T121|vTD
35806259|T121|low-dose velcade (Bortezomib), Thalidomide, Dexamethasone
35806260|T121|RVD
35806260|T121|VDR
35806260|T121|VRD
35806260|T121|VRd
35806260|T121|Revlimid (Lenalidomide), Velcade (Bortezomib), Dexamethasone
35806260|T121|Velcade (Bortezomib), Dexamethasone, Revlimid (Lenalidomide)
35806260|T121|Velcade (Bortezomib), Revlimid (Lenalidomide), Dexamethasone
35806260|T121|Velcade (Bortezomib), Revlimid (Lenalidomide), low-dose dexamethasone
35806261|T121|RVDC
35806261|T121|VDCR
35806261|T121|Revlimid (Lenalidomide), Velcade (Bortezomib), Dexamethasone, Cyclophosphamide
35806261|T121|Velcade (Bortezomib), Dexamethasone, Cyclophosphamide, Revlimid (Lenalidomide)
35806262|T121|Bisphosphonates
35806263|T121|DCEP
35806263|T121|Dexamethasone, Cyclophosphamide, Etoposide, Platinol (Cisplatin)
35806264|T121|VAD
35806264|T121|VAd
35806264|T121|Vincristine, Adriamycin (Doxorubicin), Dexamethasone
35806264|T121|Vincristine, Adriamycin (Doxorubicin), low-dose dexamethasone
35806265|T121|KTD
35806265|T121|Kyprolis (Carfilzomib), Thalidomide, Dexamethasone
35806265|T121|KTd
35806266|T121|VBMCP/VBAD
35806266|T121|Vincristine, BiCNU (Carmustine), Melphalan, Cyclophosphamide, Prednisone alternating with Vincristine, BiCNU (Carmustine), Adriamycin (Doxorubicin), Dexamethasone
35806267|T121|CVAD
35806267|T121|Cyclophosphamide, Vincristine, Adriamycin (Doxorubicin), Dexamethasone
35806268|T121|Thalidomide and Dexamethasone (TD)
35806268|T121|TD
35806268|T121|Thal-Dex
35806268|T121|Thalidomide and Dexamethasone
35806268|T121|Thalidomide, Dexamethasone
35806269|T121|PAD
35806269|T121|PAd
35806269|T121|BDD
35806269|T121|PS-341 (Bortezomib), Adriamycin (Doxorubicin), Dexamethasone
35806269|T121|PS-341 (Bortezomib), Adriamycin (Doxorubicin), low-dose dexamethasone
35806269|T121|Velcade (Bortezomib), Adriamycin (Doxorubicin), Dexamethasone
35806269|T121|Bortezomib, Doxorubicin, Dexamethasone
35806270|T121|Interferon alfa and Dexamethasone
35806271|T121|Thalidomide monotherapy
35806272|T121|VT
35806272|T121|TV
35806272|T121|Velcade (Bortezomib) and Thalidomide
35806272|T121|Thalidomide and Velcade (Bortezomib)
35806273|T121|MPR
35806273|T121|Melphalan, Prednisone, Revlimid (Lenalidomide)
35806273|T121|Melphalan, Prednisone, Lenalidomide
35806274|T121|Lenalidomide and Prednisone (RP)
35806274|T121|Revlimid (Lenalidomide) and Prednisone
35806275|T121|Tandem melphalan
35806276|T121|Antibacterials
35806277|T121|PAD (PLD substituted)
35806278|T121|EDAP
35806278|T121|Etoposide, Dexamethasone, Ara-C (Cytarabine), Platinol (Cisplatin)
35806279|T121|Bortezomib and Prednisone (VP)
35806279|T121|VP
35806279|T121|Velcade (Bortezomib) and Prednisone
35806280|T121|Carfilzomib monotherapy
35806281|T121|KCD
35806281|T121|CCyd
35806281|T121|KCyd
35806281|T121|Kyprolis (Carfilzomib), Cyclophosphamide, Dexamethasone
35806281|T121|Carfilzomib, Cyclophosphamide, dexamethasone
35806281|T121|Kyprolis (Carfilzomib), Cyclophosphamide, dexamethasone
35806282|T121|Dara-VMP
35806282|T121|D-VMP
35806282|T121|Daratumumab, Velcade (Bortezomib), Melphalan, Prednisone
35806283|T121|IRd
35806283|T121|Ixazomib, Revlimid (Lenalidomide), low-dose dexamethasone
35806284|T121|KRd
35806284|T121|Kyprolis (Carfilzomib), Revlimid (Lenalidomide), low-dose dexamethasone
35806284|T121|Carfilzomib, Revlimid (Lenalidomide), low-dose dexamethasone
35806285|T121|CPR
35806285|T121|Cyclophosphamide, Prednisone, Revlimid (Lenalidomide)
35806285|T121|REP
35806285|T121|Revlimid (Lenalidomide), Endoxan (Cyclophosphamide), Prednisone
912102|T121|Kineret
35806286|T121|MPT
35806286|T121|Melphalan, Prednisone, Thalidomide
35806287|T121|Thalidomide and Prednisolone
35806288|T121|Thalidomide and Prednisone
35806289|T121|BBD
35806289|T121|Bendamustine, Bortezomib, Dexamethasone
35806290|T121|VTP
35806290|T121|Velcade (Bortezomib), Thalidomide, Prednisone
35806291|T121|VMPT
35806291|T121|Velcade (Bortezomib), Melphalan, Prednisone, Thalidomide
912103|T121|PM-01183
912103|T121|Lurbinectedin
912104|T121|Lurbinectedin monotherapy
35806292|T121|Cyclophosphamide and G-CSF
35101743|T121|Berlex
35101742|T121|Berlocid
35806293|T121|TAD (Thalidomide)
35806293|T121|Thalidomide, Adriamycin (Doxorubicin), Dexamethasone
35806294|T121|CAD and G-CSF
35806294|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Dexamethasone
912105|T121|Metronidazole
912106|T121|Metronidazole, Tetracycline, PPI, Bismuth
35806295|T121|TVAD (Pegylated liposomal doxorubicin substituted)
35806295|T121|TVAD doxil
35806295|T121|Thalidomide, Vincristine, pegylated liposomal Adriamycin (Doxil), Dexamethasone
35806296|T121|VAD (Pegylated liposomal doxorubicin substituted)
35806296|T121|DVD
35806296|T121|DVd
35806296|T121|Doxil (Pegylated liposomal doxorubicin), Vincristine, Dexamethasone
35806296|T121|Doxil (Pegylated liposomal doxorubicin), Vincristine, low-dose dexamethasone
35806296|T121|Vincristine, Pegylated liposomal Adriamycin (Doxil), Dexamethasone
35806297|T121|VAD-P
35806297|T121|Vincristine, Adriamycin (Doxorubicin), Dexamethasone, Prednisone
35806298|T121|VAD-P/Q
35806298|T121|Vincristine, Adriamycin (Doxorubicin), Dexamethasone, Prednisone, Quinine
912107|T121|Naxitamab monotherapy
912108|T121|naxitamab-gqgk
912108|T121|Naxitamab
35806299|T121|VMP, then Rd
35806299|T121|Velcade (Bortezomib), Melphalan, Prednisone, followed by Revlimid (Lenalidomide), low dose dexamethasone
35806300|T121|VMP/Rd
35806300|T121|Velcade (Bortezomib), Melphalan, Prednisone alternating with Revlimid (Lenalidomide), low dose dexamethasone
35806301|T121|Zoledronic acid therapy
35806302|T121|BiRd
35806302|T121|C-Rd
35806302|T121|Biaxin (Clarithromycin), Revlimid (Lenalidomide), low-dose dexamethasone
35806302|T121|Clarithromycin, Revlimid (Lenalidomide), low-dose dexamethasone
35806303|T121|CYKLONE
35806303|T121|Cyclophosphamide, Kyprolis (Carfilzomib), ThaLidomide, DexamethasONE
35802851|T121|KMP
35802851|T121|CMP
35802851|T121|Kyprolis (Carfilzomib), Melphalan, Prednisone
35802851|T121|Carfilzomib, Melphalan, Prednisone
35806304|T121|Total Therapy
35806305|T121|VTD-PACE
35806305|T121|Velcade (Bortezomib), Thalidomide, Dexamethasone, Platinum (Cisplatin), Adriamycin (Doxorubicin), Cyclophosphamide, Etoposide
35101741|T121|Berofor
35806306|T121|Bortezomib and Dexamethasone (VD) and Panobinostat
35806307|T121|Bortezomib and Pegylated liposomal doxorubicin
35806308|T121|Bortezomib and Vorinostat
35806309|T121|Carfilzomib and Dexamethasone (KD)
35806310|T121|Cyclophosphamide and Dexamethasone
35806311|T121|Dara-Rd
35806311|T121|DRd
35806311|T121|Daratumumab, Revlimid (Lenalidomide), Dexamethasone
35806311|T121|D-Rd
35806311|T121|Daratumumab, Revlimid (Lenalidomide), low-dose dexamethasone
35806312|T121|Dara-VD
35806313|T121|Elo-PD
35806314|T121|Elo-Rd
35806314|T121|ELd
35806314|T121|Elotuzumab, Revlimid (Lenalidomide), low-dose dexamethasone
35806314|T121|Elotuzumab, Lenalidomide, low-dose dexamethasone
35806315|T121|Elo-VD
912109|T121|Pegfilgrastim-bmez
35806316|T121|PCD
35806316|T121|PomCyDex
35806316|T121|Pomalidomide, Cyclophosphamide, Dexamethasone
35806317|T121|Pomalidomide monotherapy
35806318|T121|Bortezomib and Cyclophosphamide
35806319|T121|BLD
35806319|T121|Bendamustine, Lenalidomide, Dexamethasone
35806320|T121|H2-receptor antagonists
35806321|T121|Bortezomib, Thalidomide, Dexamethasone, Panobinostat
35806322|T121|BTD
35806322|T121|Bendamustine, Thalidomide, Dexamethasone
35806323|T121|Carfilzomib and Panobinostat
35806324|T121|KPD
35806324|T121|CPD
35806324|T121|Kyprolis (Carfilzomib), Pomalidomide, Dexamethasone
35806324|T121|Carfilzomib, Pomalidomide, Dexamethasone
35806325|T121|CRD
35806325|T121|Cyclophosphamide, Revlimid (Lenalidomide), Dexamethasone
35806326|T121|Dara-PD
35806327|T121|DTPACE
35806327|T121|Dexamethasone, Thalidomide, Platinol (Cisplatin), Adriamycin (Doxorubicin), Cyclophosphamide, Etoposide
35806328|T121|FRD
35806328|T121|Farydak (Panobinostat), Revlimid (Lenalidomide), Dexamethasone
35806329|T121|Hyper-CVAD
35806329|T121|Hyperfractionated Cyclophosphamide, Vincristine, Adriamycin (Doxorubicin), Dexamethasone
35806330|T121|PCP
35806330|T121|Pomalidomide, Cyclophosphamide, Prednisone
35806331|T121|Pomalidomide and Prednisone
35806332|T121|PVD
35806332|T121|Pomalidomide, Velcade (Bortezomib), Dexamethasone
35806333|T121|V-HyperCAD
35806333|T121|Velcade (Bortezomib), Hyperfractionated Cyclophosphamide, Adriamycin (Doxorubicin), Dexamethasone
35806334|T121|ZRd
35806334|T121|Zolinza (Vorinostat), Revlimid (Lenalidomide), low-dose dexamethasone
35806335|T121|ABCM
35806335|T121|Adriamycin (Doxorubicin), BCNU (Carmustine), Cyclophosphamide, Melphalan
35806336|T121|mCOP/MP
35806336|T121|modified Cyclophosphamide, Oncovin (Vincristine), Prednisolone alternating with Melphalan and Prednisolone
912110|T121|Stemgen
35806337|T121|C-VAMP
35806337|T121|Cyclophosphamide, Vincristine, Adriamycin (Doxorubicin), MethylPrednisolone
35101740|T121|Bestofens
35806338|T121|DEX-IFN
35101739|T121|Bethaprim
35806339|T121|VBMCP
35806339|T121|VBCMP
35806339|T121|Vincristine, BiCNU (Carmustine), Melphalan, Cyclophosphamide, Prednisone
35806339|T121|Vincristine, BiCNU (Carmustine), Cyclophosphamide, Melphalan, Prednisone
35806340|T121|DCEP and G-CSF
35806340|T121|Dexamethasone, Cyclophosphamide, Etoposide, Platinol (Cisplatin), Granulocyte Colony Stimulating Factor
912111|T121|Tetracycline
35806341|T121|VAMP
35806341|T121|Vincristine, Adriamycin (Doxorubicin), MethylPrednisolone
35101738|T121|Bevacizumab-bvzr
35806342|T121|VBMC
35806342|T121|Vincristine, BiCNU (Carmustine), Melphalan, Cyclophosphamide
912112|T121|Tripotassium dicitratobismuthate
912113|T121|Triptorelin and RT
35806343|T121|VCP
35806344|T121|VMCP
35806344|T121|VCMP
35806344|T121|Vincristine, Melphalan, Cyclophosphamide, Prednisone
35806344|T121|Vincristine, Cyclophosphamide, Melphalan, Prednisone
35806345|T121|VMCP/VBAP
35806345|T121|Vincristine, Melphalan, Cyclophosphamide, Prednisone alternating with Vincristine, BiCNU (Carmustine), Adriamycin (Doxorubicin), Prednisone
35806346|T121|VMCP/VCAP
35806346|T121|Vincristine, Melphalan, Cyclophosphamide, Prednisone alternating with Vincristine, Cyclophosphamide, Adriamycin (Doxorubicin), Prednisone
912114|T121|UGN-101 (mitomycin-containing reverse thermal gel) monotherapy
912115|T121|Upper tract urothelial carcinoma
35806347|T121|Melphalan, then Melphalan and Busulfan
35806348|T121|MEL200, then MEL220 and Dexamethasone
35806349|T121|Melphalan, then Melphalan and TBI
35101737|T121|Bexine
35806350|T121|Melphalan, then TBI, then allo HSCT
35806351|T121|Melphalan and Methylprednisolone
35101736|T121|Beyonas Dexa
35806352|T121|Interferon alfa-2b and Prednisone
35806353|T121|Interferon alfa-2b and Thalidomide
35806354|T121|Carmustine and Doxorubicin
35806355|T121|Pomalidomide, Dexamethasone, Pembrolizumab
912116|T121|Zepzelca
35806356|T121|VAD and Cyclosporine
35806356|T121|Vincristine, Adriamycin (Doxorubicin), Dexamethasone, Cyclosporine
912117|T121|Ziextenzo
35806357|T121|CellCept
35806358|T121|ATG (Horse) monotherapy
35806358|T121|ATG
35806358|T121|AntiThymocyte Globulin
35806359|T121|ATG (Rabbit) monotherapy
35806359|T121|ATG
35806359|T121|AntiThymocyte Globulin
35806360|T121|Antibiotics
35806361|T121|Erythropoetin and Lenalidomide
35806362|T121|Busulfan and Cyclophosphamide, then allo HSCT
35101735|T121|Bibakrim
35806363|T121|DDGP
35806363|T121|Dexamethasone, DDP (Cisplatin), Gemcitabine, Pegaspargase
35806364|T121|Larotrectinib monotherapy
42542285|T121|NTRK-mutated malignancy
35806365|T121|Cesamet
35806366|T121|Fraxiparine
35806367|T121|Fraxodi
35101734|T121|Bicotrim
35806368|T121|Oxaliplatin and RT
35806368|T121|Oxaliplatin and Radiation Therapy
35806369|T121|Portrazza
35806370|T121|Aqupla
35806371|T121|Arranon
35806372|T121|Atriance
35806373|T121|Nerlynx
35806374|T121|Akynzeo
35806375|T121|GM-CSF, IL-2, Isotretinoin, Dinutuximab
35806376|T121|Isotretinoin monotherapy
35101733|T121|Bifemelan
35806377|T121|Cyclophosphamide and Vincristine
35101732|T121|Bifosa
35806378|T121|Irinotecan, Temozolomide, Dinutuximab
35101731|T121|Bifosmac
35806379|T121|Everolimus and Octreotide
35806380|T121|Fluorouracil and Streptozocin
42542286|T121|Cisplatin and Fluorouracil (CF) and Vincristine
35806381|T121|Lanreotide and Interferon alfa-2b
35806382|T121|Lanreotide monotherapy
35806383|T121|Lutetium Lu 177 dotatate and Octreotide LAR
35806383|T121|"<table class=""wikitable"" style=""color:white; background-color:#404040"">"
35806384|T121|Octreotide monotherapy
35806385|T121|Octreotide LAR monotherapy
35806386|T121|Octreotide and Interferon alfa
35806387|T121|Tasigna
35806388|T121|Anandron
35806389|T121|Nilandron
35806390|T121|Zandron
35806391|T121|Zejula
35806392|T121|Opdivo
35806393|T121|Lobectomy
35806394|T121|Pneumonectomy
35806395|T121|Lung cancer surgery
35806396|T121|Cisplatin and Vinblastine
35806396|T121|VP
35806396|T121|Vinblastine and Platinol (Cisplatin)
35806397|T121|Cisplatin and Vindesine
35806397|T121|VP
35806397|T121|VdsC
35806397|T121|Vindesine and Platinol (Cisplatin)
35806397|T121|Vindesine and Cisplatin
35806398|T121|Carboplatin, Vinorelbine, RT
35806399|T121|Cisplatin, Vinblastine, RT
35101730|T121|Bimatrim
35806400|T121|Carboplatin and Etoposide (CE)
35806400|T121|Etoposide, Paraplatin (Carboplatin)
35806400|T121|CE
35806400|T121|EC
35806400|T121|Ca/E
35806400|T121|Carboplatin and Etoposide
35806400|T121|Etoposide and Paraplatin (Carboplatin)
35806400|T121|Etoposide and Carboplatin
35806400|T121|TI-CE
35806400|T121|Taxol (Paclitaxel), Ifosfamide, Carboplatin, Etoposide
35101729|T121|Binosto
35101728|T121|Biogamma
35101727|T121|Bioprim
35101726|T121|Biosulten
35101725|T121|Biotran
35101724|T121|Biotrim
35101723|T121|Biotrin
35101722|T121|Biovorin
35101721|T121|Biprim
35806401|T121|Carboplatin and Paclitaxel (CP) and Bevacizumab
35806401|T121|Carboplatin, Paclitaxel, Bevacizumab
35806401|T121|PacCBev
35806401|T121|B+CP
35806401|T121|BCP
35806401|T121|CbTB
35806401|T121|Paclitaxel, Carboplatin, Bevacizumab
35806401|T121|Bevacizumab, Carboplatin, Paclitaxel
35806401|T121|Carboplatin, Taxol (Paclitaxel), Bevacizumab
35806401|T121|TC-BEV
35806401|T121|Taxol (Paclitaxel), Carboplatin, BEVacizumab
35806402|T121|Carboplatin and Paclitaxel (CP) and Ipilimumab
35806403|T121|Carboplatin, Pemetrexed, Pembrolizumab
35806404|T121|Pemetrexed and Pembrolizumab
35806405|T121|Carboplatin and Vinorelbine
35806405|T121|VC
35806405|T121|Vinorelbine and Carboplatin
35101720|T121|Bisbon
35101719|T121|Biseptin
35101718|T121|Biseptol
35101717|T121|Biseptrim
35101716|T121|Bismoral
35101715|T121|Bisultrim
35101714|T121|Bisuo DS
35101666|T121|Bitrim
35806406|T121|Cisplatin, Vinorelbine, Cetuximab
35806407|T121|ABCP
35806407|T121|Atezolizumab, Bevacizumab, Carboplatin, Paclitaxel
35806408|T121|Atezolizumab and Bevacizumab
35806409|T121|Carboplatin, Pemetrexed, Bevacizumab
35806409|T121|PemCBev
35806409|T121|BevCPem
35806409|T121|Pemetrexed, Carboplatin, Bevacizumab
35806409|T121|Bevacizumab, Carboplatin, Pemetrexed
35806410|T121|Pemetrexed and Bevacizumab
35806411|T121|Cisplatin and Gemcitabine (GC) and Bevacizumab
35806411|T121|GCB
35806411|T121|Gemcitabine, Cisplatin, Bevacizumab
35806412|T121|Cisplatin, Pemetrexed, Pembrolizumab
35806413|T121|Gefitinib monotherapy
35806414|T121|Carboplatin, nab-Paclitaxel, Pembrolizumab
35806415|T121|Carboplatin and Paclitaxel (CP) and Pembrolizumab
35806416|T121|Cisplatin and Gemcitabine (GC) and Necitumumab
35806417|T121|Necitumumab monotherapy
35806418|T121|Docetaxel and Nedaplatin
35806419|T121|Afatinib and Paclitaxel
35806420|T121|Amrubicin monotherapy
35806421|T121|Cabozantinib and Erlotinib
35806422|T121|Docetaxel and Vandetanib
42542287|T121|Condition
42542288|T121|ALK-positive Non-small cell lung cancer
35806423|T121|Brigatinib monotherapy
35806424|T121|Crizotinib monotherapy
35806425|T121|Lorlatinib monotherapy
42542289|T121|BRAF-mutated Non-small cell lung cancer
42542290|T121|EGFR-mutated Non-small cell lung cancer
35806426|T121|Carboplatin and Gemcitabine/Erlotinib
35806427|T121|Cisplatin and Gemcitabine/Erlotinib
35806428|T121|Dacomitinib monotherapy
35806429|T121|Gefitinib and Pemetrexed
35806429|T121|P+G
35806429|T121|Pemetrexed and Gefitinib
42542291|T121|ROS1-positive Non-small cell lung cancer
35806430|T121|MIC
35806430|T121|Mitomycin, Ifosfamide, Cisplatin
35806430|T121|Mitomycin, Ifosfamide, Platinol (Cisplatin)
35806431|T121|PEV
35806431|T121|Platinol (Cisplatin), Etoposide, Vinblastine
35806432|T121|MVP and RT
35806432|T121|Mitomycin, Vindesine, Platinol (Cisplatin), Radiation Therapy
35806433|T121|CAMP
35806433|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Methotrexate, Procarbazine
35806434|T121|CAP (Platinol)
35806434|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Platinol (Cisplatin)
35806434|T121|DCP
35806434|T121|Doxorubicin, Cyclophosphamide, Platinol (Cisplatin)
35806434|T121|Platinol (Cisplatin), Adriamycin (Doxorubicin), Cyclophosphamide
35806435|T121|Ifosfamide and Gemcitabine
35806435|T121|IG
35806436|T121|GIP
35806436|T121|Gemcitabine, Ifosfamide, Platinol (Cisplatin)
35806437|T121|MACC
35806437|T121|Methotrexate, Adriamycin (Doxorubicin), Cyclophosphamide, CCNU (Lomustine)
35101665|T121|Blexon
35806438|T121|MVP (Vinblastine)
35806438|T121|Mitomycin, Vinblastine, Platinol (Cisplatin)
35806439|T121|MVP (Vindesine)
35806439|T121|PVM
35806439|T121|Mitomycin, Vindesine, Platinol (Cisplatin)
35806439|T121|Platinol (Cisplatin), Vindesine, Mitomycin
35101664|T121|Blindafe
35806440|T121|Vindesine monotherapy
35806441|T121|VIP
35806441|T121|Vinblastine, Ifosfamide, Platinol (Cisplatin)
35806441|T121|Vepesid (Etoposide), Ifosfamide, Platinol (Cisplatin)
35806441|T121|Platinol (Cisplatin), Etoposide, Ifosfamide
35806442|T121|CR rate at 18 mo
35806443|T121|Gazyva
35806444|T121|Longastatina
35806445|T121|Octrestatin
35806446|T121|Octride
35806447|T121|Okeron
35806448|T121|Proclose
35806449|T121|Samilstin
35806450|T121|Sandostatin
35806451|T121|Sandostatina
35806452|T121|Sandostatine
35806453|T121|Longastatina LAR
35806454|T121|Sandostatin LAR
35806455|T121|Sandostatin LAR Depot
35806456|T121|Sandostatina LAR
35806457|T121|Sandostatine LAR
35806458|T121|Arzerra
35806459|T121|Zyprexa
35806460|T121|Lynparza
35806461|T121|Lartruvo
35806462|T121|Omapro
35806463|T121|Synribo
35806464|T121|Prilosec
35806465|T121|Tagrisso
35806466|T121|Cisplatin, Epirubicin, Ifosfamide
35806467|T121|MA
35806467|T121|High-dose Methotrexate, Adriamycin (Doxorubicin)
35806468|T121|MA-BCD
35806468|T121|High-dose Methotrexate, Adriamycin (Doxorubicin), Bleomycin, Cyclophosphamide, Dactinomycin
35806469|T121|MAP
35806469|T121|High-dose Methotrexate, Adriamycin (Doxorubicin), Platinol (Cisplatin)
35806470|T121|MAPIE
35806470|T121|High-dose Methotrexate, Adriamycin (Doxorubicin), Platinol (Cisplatin), Ifosfamide, Etoposide
35806471|T121|IP-BCD
35806471|T121|Ifosfamide, Platinol (Cisplatin), Bleomycin, Cyclophosphamide, Dactinomycin
35806472|T121|MAPI
35806472|T121|High-dose Methotrexate, Adriamycin (Doxorubicin), Platinol (Cisplatin), Ifosfamide
35806473|T121|M-BCD
35806473|T121|High-dose Methotrexate, Bleomycin, Cyclophosphamide, Dactinomycin
35806474|T121|M-EI
35806474|T121|Methotrexate, Etoposide, Ifosfamide
35806475|T121|MA-BCD/AP
35806475|T121|High-dose Methotrexate, Adriamycin (Doxorubicin), Bleomycin, Cyclophosphamide, Dactinomycin alternating with Adriamycin (Doxorubicin) and Platinol (Cisplatin)
35806476|T121|Cyclophosphamide and Etoposide
35806477|T121|Samarium-153 with stem cell support
35806478|T121|Ovarian cancer surgery
35806479|T121|Primary debulking surgery
35806480|T121|Altretamine monotherapy
35806481|T121|Phenothiazines
35806482|T121|Carboplatin and Gemcitabine (GCb) and Bevacizumab
35806483|T121|Carboplatin and Paclitaxel (CP) and Olaparib
35806483|T121|CP and Olaparib
35806483|T121|Carboplatin, Paclitaxel, Olaparib
35806484|T121|Rucaparib monotherapy
35806484|T121|"<table class=""wikitable"" style=""color:white; background-color:#9e4244"">"
35806485|T121|Niraparib monotherapy
35806485|T121|"<table class=""wikitable"" style=""color:white; background-color:#9e4244"">"
35806486|T121|Gemcitabine and Pegylated liposomal doxorubicin
35806487|T121|Pegylated liposomal doxorubicin and Trabectedin
35806488|T121|Paclitaxel and Pazopanib
35806489|T121|Topotecan and Bevacizumab
35806490|T121|Trabectedin monotherapy
35806491|T121|Treosulfan monotherapy
35806492|T121|Cisplatin and Cyclophosphamide
35806492|T121|CP
35806492|T121|PC
35806492|T121|Cyclophosphamide and Platinol (Cisplatin)
35806492|T121|Platinol (Cisplatin) and Cyclophosphamide
35806492|T121|CPC
35806492|T121|CisPlatin and Cyclophosphamide
35806493|T121|CHAD
35806493|T121|Cyclophosphamide, Hexalen (Altretamine), Adriamycin (Doxorubicin), DDP (Cisplatin)
35806494|T121|Chlorambucil and Cisplatin
35806495|T121|Cisplatin, Cyclophosphamide, Interferon gamma-1b
35806496|T121|Hexa-CAF
35806496|T121|Hexalen (Altretamine), Cyclophosphamide, Adrucil (Fluorouracil), Folex (Methotrexate)
35806497|T121|Altretamine and Cisplatin
912118|T121|A-CHOP
912118|T121|CHOP-C
912118|T121|Alemtuzumab, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
912118|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne, ALemtuzumab
912118|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne, Campath (Alemtuzumab)
35806498|T121|Coxatin
35806499|T121|Curaplat
35806500|T121|Cure-X
35806501|T121|Dacotin
35806502|T121|Dacplat
35806503|T121|Eloplat
35806504|T121|Eloxatin
35806505|T121|Eloxatine
35806506|T121|Oplatin
35806507|T121|OxaLitin
35806508|T121|Oxiplat
35806509|T121|Oxitan
35806510|T121|Oxzucia
35806511|T121|Sibatin
35806512|T121|Xaloplat
35806513|T121|Xylotin
35806514|T121|X-Plat
35806515|T121|Zildox
35806516|T121|Abraxane
35806517|T121|Abitaxel
35806518|T121|Altaxel
35806519|T121|Anzatax
35806520|T121|Anzatec
35806521|T121|Asotax
35806522|T121|Betaxel
35806523|T121|Bristaxol
35806524|T121|Britaxol
35806525|T121|Clitaxel
35806526|T121|Cytax
35806527|T121|Daburex
35806528|T121|Dalys
35806529|T121|Drifen
35806530|T121|Ebetaxel
35806531|T121|Formoxol
35806532|T121|Genexol
35806533|T121|Genetaxyl
35806534|T121|Gros
35806535|T121|Ifaxol
35806536|T121|Intaxel
35806537|T121|Magytax
35806538|T121|Medixel
35806539|T121|Mitotax
35806540|T121|Neotacs
35806541|T121|Neotaxan
35806542|T121|Neotaxl
35806543|T121|Ofoxel
35806544|T121|Oncotaxel
35806545|T121|Onxol
35806546|T121|Paclitax
35806547|T121|Paclitaxin
35806548|T121|Pacliteva
35806549|T121|Pacxel
35806550|T121|Padexol
35806551|T121|Paklitaxfil
35806552|T121|Panataxel
35806553|T121|Parexel
35806554|T121|Paxene
35806555|T121|Paxenor
35806556|T121|Paxus
35806557|T121|Petaxel
35806558|T121|Phyxol
35806559|T121|Poltaxel
35806560|T121|Praxel
35806561|T121|Ribotax
35806562|T121|Sindaxel
35806563|T121|Taclipaxol
35806564|T121|Tarvexol
35806565|T121|Taxocris
35806566|T121|Taxodiol
35806567|T121|Taxol
35806568|T121|Taxomedac
35806569|T121|Taycovit
35806570|T121|Unitaxel
35806571|T121|Yewtaxan
35806572|T121|Ibrance
35806573|T121|Aloxi
35806574|T121|Aredia
35806575|T121|Padium
35806576|T121|Pamisol
35806577|T121|Capecitabine and Temozolomide
35806578|T121|Doxorubicin and Streptozocin
912119|T121|Abilify
35806579|T121|FAS
35806579|T121|Fluorouracil, Adriamycin (Doxorubicin), Streptozocin
35806580|T121|Lanreotide Depot/Autogel monotherapy
912120|T121|MK-1775
912120|T121|AZD-1775
912120|T121|Adavosertib
35806581|T121|Temozolomide and Thalidomide
912121|T121|Alecinix
35806582|T121|Pancreatic cancer surgery
912122|T121|Alecnib
35806583|T121|Fluorouracil/Fluorouracil and RT
35806583|T121|Fluorouracil alternating with Fluorouracil and Radiation Therapy
35806584|T121|mFOLFIRINOX
35806584|T121|modified FOLinic acid, Fluorouracil, IRINotecan, OXaliplatin
912123|T121|Anthracenedione
35806585|T121|Gemcitabine/Fluorouracil and RT
35806585|T121|Gemcitabine alternating with Fluorouracil and Radiation Therapy
35806586|T121|Docetaxel, Gemcitabine, RT
35806586|T121|DG and RT
35806586|T121|Docetaxel, Gemcitabine, Radiation Therapy
35806587|T121|Gemcitabine, Cetuximab, RT
35806587|T121|Gemcitabine, Cetuximab, Radiation Therapy
35807526|T121|FOLFIRINOX/modified FOLFIRINOX  plus /- Chemoradiation
35807526|T121|modified FOLinic acid, Fluorouracil, IRINotecan, OXaliplatin
35806589|T121|mFOLFIRINOX, Gemcitabine, RT
35806589|T121|modified FOLinic acid, Fluorouracil, IRINotecan, OXaliplatin, Gemcitabine, Radiation Therapy
35806590|T121|Erlotinib and Gemcitabine
35806591|T121|FLEC
35806591|T121|Fluorouracil, Leucovorin (Folinic acid), Epirubicin, Carboplatin
912124|T121|Azel
912125|T121|Bdenza
912126|T121|Biganib
35101663|T121|Bolend
912127|T121|Briganix
912128|T121|Cabometyx
912129|T121|Caboxen
912130|T121|Cabozanib
912131|T121|Cabozanix
912132|T121|Cabozantinib and Nivolumab
912133|T121|CapIriRT
912133|T121|Capecitabine, Irinotecan, Radiation Therapy
912134|T121|Capmide
912135|T121|Carfilnat
912136|T121|CDK4 inhibitor
912137|T121|CDK6 inhibitor
912138|T121|Cisplatin and Fluorouracil (CF) and Pembrolizumab
912138|T121|CF and Pembrolizumab
35101661|T121|Bonaid
35101660|T121|Bonalon
35101659|T121|Bonamax
35806592|T121|GTX
35806592|T121|Gemcitabine, Taxotere (Docetaxel), Xeloda (Capecitabine)
35806593|T121|PEFG
35806593|T121|Platinol (Cisplatin), Epirubicin, Fluorouracil, Gemcitabine
42542292|T121|Docetaxel and Vinorelbine
35806594|T121|Capecitabine and Erlotinib
35101662|T121|Bonapex
35806595|T121|FULV and nanoliposomal Irinotecan
35806595|T121|5-FU, LeucoVorin (Folinic acid), nanoliposomal Irinotecan
35806596|T121|FOLFOX
35806596|T121|FOLinic acid, Fluorouracil, OXaliplatin
35806597|T121|Vectibix
35806598|T121|Faridak
35806599|T121|Farydak
35806600|T121|Protonix
35806601|T121|Votrient
35806602|T121|Oncaspar
35806603|T121|Fulphila
35806604|T121|Neulasta
35806605|T121|Onpro
35806606|T121|Pegasys
35806607|T121|PEG-Intron
35806608|T121|PegIntron
35806609|T121|Sylatron
35806610|T121|ViraferonPeg
35806611|T121|Caelyx
35806612|T121|Doxil
35806613|T121|Keytruda
35806614|T121|Alimta
35806615|T121|Antifol
35806616|T121|Kabipem
35806617|T121|Pemetero
35806618|T121|Pemetra
35806619|T121|Pemetrex
35806620|T121|Pemex
35806621|T121|Pemgem
35806622|T121|Pemibenz
35806623|T121|Pemnat
35806624|T121|Pexotra
35806625|T121|TIP
35806625|T121|Taxol (Paclitaxel), Ifosfamide, Platinol (Cisplatin)
35806626|T121|VBM (Vincristine)
35806626|T121|VBM
35806626|T121|Vincristine, Bleomycin, Methotrexate
35806627|T121|BMP
35806627|T121|MPB
35806627|T121|Bleomycin, Methotrexate, Platinol (Cisplatin)
35806627|T121|Methotrexate, Platinol (Cisplatin), Bleomycin
35806628|T121|Benambax
35806629|T121|Lomidine
35806630|T121|Nebupent
35806631|T121|Pentam
35806632|T121|Pentamidina
35806633|T121|Pneumopent
35806634|T121|Nipent
35101658|T121|Bonemax
35806635|T121|CMED
35806635|T121|Cyclophosphamide, Methotrexate, Etoposide, Dexamethasone
35806636|T121|GDPT
35806636|T121|Gemcitabine, DDP (Cisplatin), Prednisone, Thalidomide
35806637|T121|CHOP and Everolimus
35806637|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne, Everolimus
35806638|T121|CHOP-AL
35806639|T121|HyperCHidam
35806639|T121|Hyperfractionated Cyclophosphamide, Hiigh-dose ara-c (Cytarabine) and methotrexate
35806640|T121|DD-CHOP
35806640|T121|Denileukin, Diftitox, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
35806588|T121|TFC, then allo HSCT
35806588|T121|TFC
35806588|T121|Thiotepa, Fludarabine, Cyclophosphamide
35806641|T121|Bortezomib and Panobinostat
35806642|T121|Chidamide monotherapy
35101657|T121|Bongard
35806643|T121|Forodesine monotherapy
912139|T121|CHOP-14 (Prednisolone)
912139|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisolone every 14 days
35806644|T121|Omnitarg
35806645|T121|Perjeta
35806646|T121|Cyclophosphamide, Dacarbazine, Vincristine
35806646|T121|CVD
35806646|T121|Cyclophosphamide, Vincristine, Dacarbazine
35806647|T121|AquaMephyton
35806648|T121|Konakion
35806649|T121|Pinorubicin
35806650|T121|Pinorubin
35806651|T121|Therarubicin
35806652|T121|Pixuvri
35806653|T121|PAD/VCD
35806653|T121|PS-341 (Bortezomib), Adriamycin liposomal (Pegylated liposomal doxorubicin), Dexamethasone alternating with Velcade (Bortezomib), Cyclophosphamide, Dexamethasone
35806654|T121|Mozobil
35806655|T121|Aspirin monotherapy
35806656|T121|Interferon monotherapy
35101656|T121|Bonmax
35806657|T121|Actimid
35806658|T121|Ibipolid
35806659|T121|Imnovid
35806660|T121|Pomalid
35806661|T121|Pomalyst
35806662|T121|Iclusig
35806663|T121|ACVBP, dose-adjusted
35806663|T121|Adriamycin (Doxorubicin), Cyclophosphamide, Vindesine, Bleomycin, Prednisone
35806664|T121|R, then CHOP
35806664|T121|Rituximab followed by Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Predniso(lo)ne
35806665|T121|R-CP
35806665|T121|Rituximab, Cyclophosphamide, Prednisone or Prednisolone
35806666|T121|Reduction of immunosuppression
35806666|T121|RIS
35806666|T121|Reduction of ImmunoSuppression
35806667|T121|Folotyn
35806668|T121|Effient
35806669|T121|Efient
35806670|T121|Glitax
35806671|T121|Prasita
35806672|T121|Prasudoc
35806673|T121|PrasuSafe
35806674|T121|Prax
35806675|T121|Surfent
35806676|T121|Targol
35806677|T121|Pravachol
35806678|T121|Adnisolone
35806679|T121|Aprednislon
35806680|T121|Capsoid
35806681|T121|Cortalone
35806682|T121|Cortisolone
35806683|T121|Cotolone
35806684|T121|Dacortin H
35806685|T121|Decaprednil
35806686|T121|Decortin H
35806687|T121|Delta-Cortef
35806688|T121|Deltacortril
35806689|T121|Delta-Diona
35806690|T121|Delta-Phoricol
35806691|T121|Deltasolone
35806692|T121|Deltidrosol
35806693|T121|Dhasolone
35806694|T121|Di-Adreson-F
35806695|T121|Dontisolon D
35806696|T121|Estilsona
35806697|T121|Fisopred
35806698|T121|Frisolona
35806699|T121|Gupisone
35806700|T121|Hostacortin H
35806701|T121|Hydeltra
35806702|T121|Hydeltrasol
35806703|T121|Klismacort
35806704|T121|Kuhlprednon
35806705|T121|Lenisolone
35806706|T121|Lepi-Cortinolo
35806707|T121|Linola-H N
35806708|T121|Linola-H-Fett N
35806709|T121|Longiprednil
35806710|T121|Medicort
35806711|T121|Meticortelone
35806712|T121|Meti-derm
35806713|T121|Millipred
35806714|T121|Opredsone
35806715|T121|Orapred
35806716|T121|Panafcortelone
35806717|T121|Predcor
35806718|T121|Predicort
35806719|T121|Precortisyl
35806720|T121|Pred-Clysma
35806721|T121|Predeltilone
35806722|T121|Predni-Coelin
35806723|T121|Prednicortelone
35806724|T121|Predni-Helvacort
35806725|T121|Prelone
35806726|T121|Prenilone
35806727|T121|Pri-Cortin
35806728|T121|Veripred
35806729|T121|Artinizona
35806730|T121|Artrizona
35806731|T121|Becortem
35806732|T121|Bersen
35806733|T121|Colisone
35806734|T121|Cortancyl
35806735|T121|Corticorten
35806736|T121|Cortigen
35806737|T121|Cortiol
35806738|T121|Cortiprex
35806739|T121|Cutason
35806740|T121|Dacortin
35806741|T121|Decortancyl
35806742|T121|Decortin
35806743|T121|Decortisyl
35806744|T121|Dehydrocortison
35806745|T121|Delcortin
35806746|T121|Dellacorta
35806747|T121|Delta-Cortisone
35806748|T121|Delta Cortelan
35806749|T121|Deltacortene
35806750|T121|Deltacortone
35806751|T121|Deltason
35806752|T121|Deltasone
35806753|T121|Deltisona
35806754|T121|Dispersona
35806755|T121|Drazone
35806756|T121|Econosone
35806757|T121|Ednaprom
35806758|T121|Encorton
35806759|T121|Erlanison
35806760|T121|Flamacorten
35806761|T121|Hostacortin
35806762|T121|Ifison
35806763|T121|Isolone
35806764|T121|Lisacort
35806765|T121|ME Korti
35806766|T121|Meticorten
35806767|T121|Nisocortec
35806768|T121|Nisona
35806769|T121|Nisone
35806770|T121|Nizon
35806771|T121|Nosipren
35806772|T121|Novoprednisone
35806773|T121|Orasone
35806774|T121|Panafcort
35806775|T121|Panasol-S
35806776|T121|Pehacort
35806777|T121|Pharmapred
35806778|T121|Precortil
35806779|T121|Predcort
35806780|T121|Predeltin
35806781|T121|Predicor
35806782|T121|Predicorten
35806783|T121|Predinis
35806784|T121|Preditec
35806785|T121|Prednax
35806786|T121|Prednicap
35806787|T121|Prednicen-M
35806788|T121|Prednilonga-Retard
35806789|T121|Predniment
35806790|T121|Prednison
35806791|T121|Prednisona
35806792|T121|Prednisonum
35806793|T121|Prednitone
35806794|T121|Predson
35806795|T121|Predsone
35806796|T121|Predval
35806797|T121|Procion
35806798|T121|Prolix
35806799|T121|Pronison
35806800|T121|Pulmison
35806801|T121|Rectodelt
35806802|T121|Senterlic
35806803|T121|Sone
35806804|T121|Steerometz
35806805|T121|Sterapred
35806806|T121|Trolic
35806807|T121|Ultracorten
35806808|T121|Vitazon
35806809|T121|Winpred
35806810|T121|Indicarb
35806811|T121|Matulane
35806812|T121|Natulan
35806813|T121|Natulanar
35806814|T121|P-Carzine
35806815|T121|Acuvert
35806816|T121|Compazine
35806817|T121|Compro
35806818|T121|Dvometil
35806819|T121|Stemetil
35806820|T121|Phenergan
35806821|T121|ADT
35806821|T121|Androgen Deprivation Therapy
35806822|T121|ADT and RT
35806822|T121|Androgen Deprivation Therapy and Radiation Therapy
35806823|T121|Flutamide and Goserelin
35806824|T121|Active surveillance
35101655|T121|Bonomax
35806825|T121|GnRH antagonists
35806826|T121|Bilateral orchiectomy
35806827|T121|Flutamide, Goserelin, RT
35806827|T121|Flutamide, Goserelin, Radiation Therapy
912140|T121|CK1 epsilon inhibitor
912141|T121|CK1 inhibitor
35806828|T121|Flutamide, Leuprolide, RT
35806828|T121|Flutamide, Leuprolide, Radiation Therapy
35806829|T121|Goserelin and RT
35806829|T121|Goserelin and Radiation Therapy
35806830|T121|Bicalutamide and Goserelin
35806831|T121|Radical prostatectomy
35806832|T121|Bicalutamide and RT
35806832|T121|Bicalutamide and Radiation Therapy
35806833|T121|Prostatectomy with lymphadenectomy
35806834|T121|Prostatectomy
35806835|T121|ADT and Apalutamide
35806835|T121|Androgen Deprivation Therapy and Apalutamide
35806836|T121|ADT and Enzalutamide
35806836|T121|Androgen Deprivation Therapy and Enzalutamide
35806837|T121|ADT and Abiraterone
35806837|T121|Androgen Deprivation Therapy and Abiraterone
35806838|T121|ADT and Docetaxel
35806838|T121|Androgen Deprivation Therapy and Docetaxel
35806839|T121|Docetaxel, Estramustine, Goserelin
35806840|T121|Bicalutamide monotherapy
35101654|T121|Benralizumab
35101653|T121|Benralizumab monotherapy
35101652|T121|Fasenra
35806841|T121|Bicalutamide and Leuprolide
35806842|T121|Degarelix monotherapy
35806843|T121|Flutamide monotherapy
35806844|T121|Flutamide and Leuprolide
912142|T121|Colchicine
35806845|T121|Intermittent ADT
35806845|T121|IHT
35806845|T121|Intermittent Hormone Therapy
35806846|T121|Nonsteroidal antiandrogens
35806847|T121|Nilutamide and Orchiectomy
912143|T121|Colcrys
35806848|T121|Abiraterone monotherapy
35806849|T121|Antiandrogen withdrawal
35806850|T121|Apalutamide monotherapy
35806851|T121|Hydrocortisone monotherapy
35806852|T121|Ketoconazole and Hydrocortisone
35806853|T121|Ketoconazole, Hydrocortisone, Dutasteride
35806854|T121|Cabazitaxel and Prednisone
35806855|T121|Carboplatin, Docetaxel, Prednisone
35101651|T121|Boschtrim
912144|T121|Cometriq
35806856|T121|Cyclophosphamide, Prednisone, Diethylstilbestrol
35806856|T121|CPD
35806857|T121|Docetaxel and Estramustine
35806858|T121|Docetaxel and Prednisone
35806859|T121|Mitoxantrone and Prednisone
35806860|T121|Ipilimumab and RT
35806860|T121|Ipilimumab and Radiation Therapy
35806861|T121|Sipuleucel-T monotherapy
35806862|T121|Radium-223 monotherapy
35806863|T121|Samarium-153 monotherapy
35101650|T121|Bostrong
35806864|T121|Aspirin and Dexamethasone
35806864|T121|DA
35806864|T121|Dexamethasone and Aspirin
35806865|T121|Castration
35806866|T121|Cortisone monotherapy
35806867|T121|Cyproterone acetate monotherapy
35806868|T121|Doxorubicin and Strontium-89
35806869|T121|Beriplex
35806870|T121|Confidex
35806871|T121|Kcentra
35806872|T121|Octaplex
35806873|T121|Profilnine
35806874|T121|Alpharadin
35806875|T121|Xofigo
35806876|T121|Supect
35806877|T121|Tomudex
35806878|T121|IBset
35806879|T121|Iribo
35806880|T121|Nasea
35806881|T121|Nozia
35806882|T121|Cyramza
35806883|T121|Cymer
35806884|T121|Cymerin
35806885|T121|Elitek
35806886|T121|Fasturtec
35806887|T121|Rasbelon
35806888|T121|Rasburnat
35806889|T121|Rasby
35806890|T121|Capecitabine and RT
35806890|T121|Capecitabine and Radiation Therapy
35806891|T121|Rectal cancer surgery
35806892|T121|Capecitabine, Sorafenib, RT
35806892|T121|Capecitabine, Sorafenib, Radiation Therapy
35806893|T121|CapeOx, Cetuximab, RT
35806893|T121|CapeOX, Cetuximab, RT
35806893|T121|Capecitabine, OXaliplatin, Cetuximab, Radiation Therapy
35806894|T121|FULV and RT
35806894|T121|FluoroUracil, LeucoVorin (Folinic acid) and Radiation Therapy
35806895|T121|mFOLFOX6 and RT
35806895|T121|modified FOLinic acid, Fluorouracil, OXaliplatin and Radiation Therapy
35806896|T121|UFT monotherapy
35806897|T121|Capecitabine/Capecitabine and RT
35806897|T121|Capecitabine alternating with Capecitabine and Radiation Therapy
35806898|T121|Fluorouracil, then Fluorouracil and RT, then Fluorouracil
35806899|T121|Renal cell carcinoma surgery
35806900|T121|Axitinib and Avelumab
35806901|T121|Axitinib monotherapy
35806902|T121|Bevacizumab and Interferon alfa-2a
35806903|T121|Doxorubicin and Gemcitabine
35806904|T121|Gemcitabine and Sunitinib
35806905|T121|Interferon alfa-2a and Interleukin-2
35806906|T121|Everolimus and Lenvatinib
35806907|T121|Interferon alfa-2a and Isotretinoin
35806908|T121|Interferon alfa-2c monotherapy
35806909|T121|VA
35806909|T121|Vincristine and Actinomycin D
35806910|T121|VAC
35806910|T121|Vincristine, Actinomycin D, Cyclophosphamide
35806911|T121|VI, then VDC/IE, then VAC, then VI
35806911|T121|Vincristine and Irinotecan, followed by Vincristine, Doxorubicin, Cyclophosphamide alternating with Ifosfamide and Etoposide, followed by Vincristine, Actinomycin D, Cyclophosphamide, followed by Vincristine and Irinotecan
35806912|T121|VIE
35806912|T121|Vincristine, Ifosfamide, Etoposide
35806913|T121|Kisqali
35806914|T121|Truxima
35806915|T121|Ikgdar
35806916|T121|Mabtas
35806917|T121|MabThera
35806918|T121|Reditux
35806919|T121|Ristova
35806920|T121|Rituxan
35806921|T121|Rituxim
35806922|T121|Transera-Kit
35806923|T121|Xarelto
35806924|T121|Varubi
35806925|T121|Varubi IV
35806926|T121|Istodax
35806927|T121|Rubraca
35806928|T121|Jakafi
35806929|T121|Jakavi
42542293|T121|Hedgehog pathway-mutated malignancy
35806930|T121|Quadramet
35806931|T121|Leukine
35806932|T121|Scopoderm
35806933|T121|Transderm Scop
35806934|T121|Semustina
35806935|T121|L-glutamine monotherapy
35806936|T121|Sylvant
35806937|T121|Provenge
35806938|T121|Rapamune
35806939|T121|CEV and RT
35806939|T121|Cyclophosphamide, Epirubicin, Vincristine, Radiation Therapy
35806940|T121|Belotecan and Cisplatin
35806940|T121|Belotecan and Platinol (Cisplatin)
35806941|T121|Carboplatin and Etoposide (CE) and Atezolizumab
35806941|T121|CE and Atezolizumab
35806941|T121|Carboplatin, Etoposide, Atezolizumab
35806942|T121|Carboplatin and Etoposide (CE) Bevacizumab
35806943|T121|Carboplatin and Irinotecan
35806943|T121|IC
35806943|T121|Irinotecan and Carboplatin
35806943|T121|Irinotecan and Paraplatin (Carboplatin)
35806944|T121|CAV
35806944|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Vincristine
35806944|T121|Vincristine, Adriamycin (Doxorubicin), Cyclophosphamide
35806944|T121| CAO
35806944|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Oncovin (Vincristine)
35101649|T121|Bendamustine and Rituximab (BR) and Polatuzumab vedotin
35101649|T121|BR and Polatuzumab vedotin
35101649|T121|Bendamustine, Rituximab, Polatuzumab vedotin
35806945|T121|Cisplatin and Etoposide (EP) and Bevacizumab
35806946|T121|Teniposide monotherapy
35806947|T121|Cisplatin, Etoposide, Irinotecan
35806948|T121|Epirubicin and Ifosfamide
35806948|T121|EI
35806948|T121|Epirubicin, Ifosfamide
912145|T121|DepoCyt
912146|T121|Diamox
35806949|T121|VMV-VAC
35806949|T121|Vincristine, Methotrexate, VP-16 (Etoposide), VP-16 (Etoposide), Adriamycin (Doxorubicin), Cyclophosphamide
35806950|T121|CC/DE and RT
35806950|T121|Cyclophosphamide and Cisplatin alternating with Doxorubicin and Etoposide, with Radiation Therapy
35806951|T121|Methotrexate, RT, Cyclophosphamide
35806952|T121|BACO
35806952|T121|Bleomycin, Adriamycin (Doxorubicin), Cyclophosphamide, Oncovin (Vincristine)
35806953|T121|CAV/PE
35806953|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Vincristine alternating with Platinol (Cisplatin) and Etoposide
35806954|T121|CDE
35806954|T121|CAE
35806954|T121|Cyclophosphamide, Doxorubicin, Etoposide
35806954|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Etoposide
35806956|T121|CEV (Cyclophosphamide/Epirubicin)
35806956|T121|CEV
35806956|T121|Cyclophosphamide, Epirubicin, Vincristine
35806957|T121|CEV (Carboplatin/Etoposide)
35806957|T121|CEV
35806957|T121|Carboplatin, Etoposide, Vincristine
35806958|T121|Cyclophosphamide, Lomustine, Methotrexate
35806959|T121|EVI
35806959|T121|Epirubicin, Vindesine, Ifosfamide
35806960|T121|PCDE
35806960|T121|Platinol (Cisplatin), Cyclophosphamide, EpiDoxorubicin (Epirubicin), Etoposide
35806961|T121|TEC
35806962|T121|EIA
35806962|T121|Etoposide, Ifosfamide, Adriamycin (Doxorubicin)
42542294|T121|FOLFOXIRI and Panitumumab
42542294|T121|FOLinic acid, Fluorouracil, OXaliplatin, IRInotecan, Panitumumab
35806964|T121|Dacarbazine and Doxorubicin
35806964|T121|AD
35806964|T121|Adriamycin (Doxorubicin) and Dacarbazine
35806965|T121|Doxorubicin and Ifosfamide
35806965|T121|Adriamycin (Doxorubicin), Ifosfamide, Mesna
35806966|T121|Doxorubicin, Ifosfamide, RT
35806966|T121|AIM and RT
35806966|T121|Adriamycin (Doxorubicin), Ifosfamide, Mesna, Radiation Therapy
35806967|T121|Doxorubicin and Olaratumab
35806968|T121|MAID
35806968|T121|Mesna, Adriamycin (Doxorubicin), Ifosfamide, Dacarbazine
35806969|T121|Dacarbazine and Gemcitabine
35806970|T121|Odomzo
35806955|T121|Nexavar
35806963|T121|Sorafenat
35806971|T121|Soranib
35806972|T121|Cytarabine, Ifosfamide, G-CSF
35806973|T121|CYVE and G-CSF
35806973|T121|CYtarabine, VEpesid (Etoposide), Granulocyte Colony Stimulating Factor
35806974|T121|IGEV and G-CSF
35806974|T121|Ifosfamide, GEmcitabine, Vinorelbine, Granulocyte Colony Stimulating Factor
35806975|T121|Zanosar
35806976|T121|Suninat
35806977|T121|Sutent
35806978|T121|Cyclophosphamide, Cytarabine, Mercaptopurine, Pegaspargase, Vincristine
35806979|T121|Cyclophosphamide, Cytarabine, Mercaptopurine, Nelarabine, Pegaspargase, Vincristine
35806980|T121|Doxorubicin, L-asparaginase, Mercaptopurine, Methotrexate, Vincristine, Prednisone
35806981|T121|L-asparaginase monotherapy
35806982|T121|Methotrexate, Pegaspargase, Vincristine
35806982|T121|COG C-MTX
35806982|T121|Children's Oncology Group Capizzi-style MTX (Methotrexate) regimen
35806983|T121|Nelarabine monotherapy
35806984|T121|Advagraf
35806985|T121|Prograf
35806986|T121|Elzonris
35806987|T121|Talzenna
35806988|T121|Imlygic
35806989|T121|OncoVEX^GM-CSF
35806990|T121|Amnoid
35806991|T121|Amnolake
35806992|T121|Istubal
35806993|T121|Nolvadex
35806994|T121|Soltamox
35806995|T121|Valodex
35806996|T121|Granix
35806997|T121|Neutroval
35806998|T121|Teysuno
35806999|T121|Ftorafur
35807000|T121|Luporal
35807001|T121|Tefudex
35807002|T121|Ufur
35807003|T121|Uftoral
35807004|T121|Uracel
35807005|T121|Xermelo
35807006|T121|Gliotem
35807007|T121|Temcad
35807008|T121|Temizole
35807009|T121|Temodal
35807010|T121|Temodar
35807011|T121|Temonat
35807012|T121|Temoside
35807013|T121|Temoz
35807014|T121|Temzol
35807015|T121|Vumon
35807016|T121|C-BOP
35807016|T121|Cisplatin, Bleomycin, Oncovin (Vincristine), Paraplatin (Carboplatin)
35807017|T121|Accelerated BEP
35807017|T121|Accelerated Bleomycin, Etoposide, Platinol (Cisplatin)
35807018|T121|Bleomycin and Vincristine (BO)
35807018|T121|BO
35807018|T121|Bleomycin and Oncovin (Vincristine)
35807019|T121|M-TIP
35807019|T121|Methotrexate, Taxol (Paclitaxel), Ifosfamide, Platinol (Cisplatin)
35101648|T121|Brek
35807020|T121|PVeBV
35807020|T121|VBEP
35807020|T121|Platinol (Cisplatin), Velban (Vinblastine), Bleomycin, Vepesid (Etoposide)
35807020|T121|Vinblastine, Bleomycin, Etoposide, Platinol (Cisplatin)
35807021|T121|Carboplatin and Etoposide, then auto HSCT
35807022|T121|Cisplatin and Epirubicin
35807022|T121|CIS-EPI
35807022|T121|CISplatin, EPIrubicin
35807023|T121|VeIP
35807023|T121|Velban (Vinblastine), Ifosfamide, Platinol (Cisplatin)
35807024|T121|Gemcitabine, Oxaliplatin, Paclitaxel
35807024|T121|GOP
35807025|T121|Oxaliplatin and Bevacizumab
35807026|T121|BVP
35807026|T121|PVB
35807026|T121|Bleomycin, Vinblastine, Platinol (Cisplatin)
35807026|T121|Platinol (Cisplatin), Vinblastine, Bleomycin
35807026|T121|Vinblastine, Bleomycin, DDP (Cisplatin)
35807027|T121|Bleomycin and Vinblastine
35807028|T121|Chlorambucil, Dactinomycin, Methotrexate
35807029|T121|CISCA/VB
35807029|T121|CISplatin, Cyclophosphamide, Adriamycin (Doxorubicin) alternating with Vinblastine and Bleomycin
35807030|T121|Plicamycin monotherapy
35807031|T121|Thaangio
35807032|T121|Thalide
35807033|T121|Thalix
35807034|T121|Thalomid
35807035|T121|Zuvimide
35807036|T121|Tabloid
35807037|T121|Tepadina
35807038|T121|Thioplex
35807039|T121|Lusutrombopag monotherapy
35807040|T121|Plasma exchange
912147|T121|Enzamide
35807041|T121|Caplacizumab and Plasma exchange
35807042|T121|Methylprednisolone monotherapy
35807043|T121|Vincristine monotherapy
35807044|T121|PAC
35807044|T121|Platinol (Cisplatin), Adriamycin (Doxorubicin), Cyclophosphamide
35807044|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Platinol (Cisplatin)
35807045|T121|Thymectomy
35807046|T121|ADOC
35807046|T121|Adriamycin (Doxorubicin), cis-Diamminedichloroplatinum (Cisplatin), Oncovin (Vincristine), Cyclophosphamide
35101647|T121|Brifeseptol
35807047|T121|Octreotide and Prednisone
35807048|T121|Radioiodine ablation
35807049|T121|Thyroidectomy
35807050|T121|Vandetanib monotherapy
42542295|T121|BRAF-mutated Thyroid cancer
35807051|T121|Ticlid
35807052|T121|Tilopin
35807053|T121|Innohep
35807054|T121|Tinprin
35807055|T121|Aggrastat
35807056|T121|Kymriah
35807057|T121|Xeljanz
35807058|T121|Acapodene
35807059|T121|Fareston
35807060|T121|Bexxar
35807061|T121|Yondelis
35807062|T121|Mekinist
35807063|T121|Herzuma
35807064|T121|Biceltis
35807065|T121|CANMab
35807066|T121|Herceptin
35807067|T121|Herclon
35807068|T121|Hertraz
35807069|T121|Ovastat
35807070|T121|Trecondi
35807071|T121|Lonsurf
35807072|T121|Decapeptyl
35807073|T121|Diphereline
35807074|T121|Gonapeptyl
35807075|T121|Trelstar LA
35807076|T121|Variopeptyl
35807077|T121|Abatoarin
35807078|T121|Hensetron
35807079|T121|Navoban
35807080|T121|Setrovel
35807081|T121|Vistogard
35807082|T121|Talavir
35807083|T121|Valcivir
35807084|T121|Valtrex
35807085|T121|Virval
35807086|T121|Zelitrex
35807087|T121|Caprelsa
35807088|T121|Zactima
35807089|T121|ABV (Vinblastine)
35807089|T121|Adriamycin (Doxorubicin), Bleomycin, Vinblastine
35807090|T121|ABV (Vincristine)
35807090|T121|Adriamycin (Doxorubicin), Bleomycin, Vincristine
35807092|T121|Daunorubicin liposomal monotherapy
35807091|T121|Zelboraf
35807093|T121|Venclexta
35807094|T121|Apixaban monotherapy
35807095|T121|Betrixaban monotherapy
35807096|T121|Enoxaparin monotherapy
35807097|T121|Dalteparin monotherapy
35807098|T121|Bivalirudin monotherapy
35807099|T121|Dabigatran monotherapy
35807100|T121|Edoxaban monotherapy
35807101|T121|Heparin monotherapy
35807101|T121|UnFractionated Heparin
35807102|T121|Tinzaparin monotherapy
35802852|T121|Alkaban-AQ
35807103|T121|Blastovin
35807104|T121|Cellblastin
35807105|T121|Cytoblastine
35807106|T121|Erbablas
35807107|T121|Exal
35807108|T121|Faulblastina
35807109|T121|Lemblastine
35807110|T121|Periblastine
35807111|T121|Rabinefil
35807112|T121|Velban
35807113|T121|Velbastine
35807114|T121|Velbe
35807115|T121|Vinblasin
35807116|T121|Vinblastin
35807117|T121|Vinblastina
35807118|T121|Alcrist
35807119|T121|Biocrist
35807120|T121|Biocrystin
35807121|T121|Cellcristin
35807122|T121|Citomid
35807123|T121|Crivosin
35807124|T121|Farmistin CS
35807125|T121|Fauldvincri
35807126|T121|Krebin
35807127|T121|Kyocristine
35807128|T121|Nevexitin
35807129|T121|Onkocristin
35807130|T121|Pericristine
35807131|T121|Pharmacristine
35807132|T121|Tecnocris
35807133|T121|Vincasar
35807134|T121|Vinces
35807135|T121|Vincosid
35807136|T121|Vincran
35807137|T121|Vincrex
35807138|T121|Vincrifil
35807139|T121|Vincrin
35807140|T121|Vincrisin
35807141|T121|Vincrisol
35807142|T121|Vincristin
35807143|T121|Vincristina
35807144|T121|Vincristinesulfaat
35807145|T121|Vincristinsulfat
35807146|T121|Vincristinum
35807147|T121|Vincrisul
35807148|T121|Vinracin
35807149|T121|Vinracine
35807150|T121|Vinstin
35807151|T121|Vintec
35807152|T121|Marqibo
35807153|T121|Eldesine
35807154|T121|Eldisin
35807155|T121|Enison
35807156|T121|Fildesin
35807157|T121|Gesidine
35807158|T121|Erivedge
35807159|T121|antihemophilic factor/von Willebrand Factor complex
35807159|T121|Von Willebrand factor and factor VIII complex human
35807160|T121|Alphanate
35807161|T121|Humate-P
35807162|T121|Wilate
35807163|T121|Wilfactin
35807164|T121|Zontivity
35807165|T121|Zolinza
35807166|T121|Plerixafor monotherapy
35807167|T121|CaRD
35807167|T121|Carfilzomib, Rituximab, Dexamethasone
35807168|T121|DRC
35807168|T121|Dexamethasone, Rituximab, Cyclophosphamide
35101646|T121|Broncoflam
35101645|T121|Brongenit
35807169|T121|Thalidomide and Rituximab
35807170|T121|Thioguanine monotherapy
912148|T121|HH-GV-678
912148|T121|flumatinib mesylate
912148|T121|Flumatinib
35807171|T121|RVR
35807171|T121|RAD-001 (Everolimus), Velcade (Bortezomib), Rituximab
35807172|T121|Dactinomycin and Vincristine
35807173|T121|Aztec
35807174|T121|Retrovir
35807175|T121|Eylea
35807176|T121|Zaltrap
35807177|T121|Aclasta
35807178|T121|Blaztere
35807179|T121|Cytozol
35807180|T121|Reclast
35807181|T121|Servycal
35807182|T121|Zobone
35807183|T121|Zoldonat
35807184|T121|Zomera
35807185|T121|Zometa
35807186|T121|Zyfoss
35101644|T121|mFOLFOX6 (L-Leucovorin)
35101644|T121|modified FOLinic acid, Fluorouracil, OXaliplatin
35101644|T121|modified L-FOLinic acid, Fluorouracil, OXaliplatin
35101643|T121|mFOLFOX6-B (L-Leucovorin)
35101643|T121|FOLFOX-B
35101643|T121|modified L-FOLinic acid, Fluorouracil, OXaliplatin, Bevacizumab
35101643|T121|FOLinic acid, Fluorouracil, OXaliplatin, Bevacizumab
35101642|T121|mFOLFOX7 (L-Leucovorin)
35101642|T121|modified L-FOLinic acid, Fluorouracil, OXaliplatin
35101641|T121|Plerixafor and G-CSF
42542296|T121|Gastroesophageal cancer
42542297|T121|Gemcitabine and S-1
42542297|T121|GS
35101640|T121|TH-FEC (Docetaxel, SC Trastuzumab)
35101640|T121|TH-FEC
35101640|T121|Taxotere (Docetaxel) and Herceptin Hylecta (Trastuzumab and hyaluronidase), followed by Fluorouracil, Epirubicin, Cyclophosphamide
35101639|T121|Trastuzumab and hyaluronidase monotherapy
42542298|T121|Allogeneic stem cells
42542299|T121|BID
42542299|T121|Bendamustine, Ixazomib, Dexamethasone
912149|T121|Carboplatin and Etoposide (CE) and Thalidomide
42542300|T121|Doxorubicin and Fluorouracil
35101638|T121|Brulin
35101637|T121|Bryterol
35101636|T121|BS
35101635|T121|Buateron
912150|T121|FUDR
35101634|T121|Bucokon
35101633|T121|131I-Metaiodobenzylguanidine (131I-MIBG)
35101632|T121|Bufadexon
912151|T121|Gastric MALT lymphoma, H. Pylori eradication therapy
35101631|T121|Butiol
35101630|T121|CA ATRA
35101629|T121|Calc Leucovorn
35101628|T121|Calcifolin
35101627|T121|Calcium Folinato
35101626|T121|Calcium Folint
35101625|T121|Calcium Leucovorin
35101624|T121|Calcium Leucovorn
35101623|T121|Calciumfolin
35101622|T121|Calciumfolinat
35101621|T121|Calcivoran
35101620|T121|Calfolex
35101619|T121|Calfolin
35101618|T121|Calidron
35101617|T121|Calinat
35101616|T121|Canalon
35101615|T121|Canferon A
35101614|T121|Canprim
912152|T121|Glenza
35101613|T121|Carbidu
35101612|T121|Carboplatin, Etoposide, RT
35101612|T121|EP and RT
35101612|T121|Etoposide, Paraplatin (Carboplatin), Radiation Therapy
35101611|T121|Carboplatin, nab-Paclitaxel, Atezolizumab
35101611|T121|A+CnP
35101611|T121|Atezolizumab, Carboplatin, nab-Paclitaxel
35101610|T121|Caretran
35101609|T121|Carulon
35101608|T121|Caumadin
912153|T121|HER2-positive Gastric cancer
35101607|T121|Cebedex
35101606|T121|Cedantron
35101605|T121|Cefixime
35101604|T121|Cehafolin
35101603|T121|Cellacort
35101602|T121|Celudex
35101601|T121|Centrim
35101600|T121|Cephalexin
35101599|T121|Cephalosporin
35101598|T121|Ceramos
35101597|T121|Cetadexon
42542301|T121|Malignant breast neoplasm
42542302|T121|Malignant solid neoplasm
35101596|T121|Chemitrim
35101595|T121|Chemix
35101594|T121|Chemizol
35101593|T121|Chemoprim
35101592|T121|Chemotran
35101591|T121|Chemotrim
35101590|T121|Chemotrin
35101589|T121|Chemozole
35807188|T121|Chemotherapeutic
35807189|T121|Immunotherapeutic
35807190|T121|Antibody medication
35807191|T121|T-cell activator
35807192|T121|BiTE antibody
35807193|T121|Anti-CD33 antibody
35807194|T121|Anti-CD3 antibody
35807195|T121|Investigational drug
35807196|T121|Oral
35807197|T121|Kinase inhibitor
35807198|T121|AKT1 inhibitor
35807199|T121|Intravenous
35807200|T121|GPIIb-IIIa inhibitor
35807201|T121|Anti-GPIIb-IIIa antibody
35807202|T121|Protein expression-specific medication
35807203|T121|CDK inhibitor
35807204|T121|HDAC inhibitor
35807205|T121|Endocrine therapeutic
35807206|T121|Antiandrogen
35807207|T121|Steroid synthesis inhibitor
35807208|T121|BTK inhibitor
35807209|T121|Rectal
35807210|T121|Antipyretic
35807211|T121|FDA approved drug
35807212|T121|OTC medication
35807213|T121|WHO Essential Pain and Palliative Care Medicine
35807214|T121|Anthracycline
35807215|T121|Topoisomerase inhibitor
35807216|T121|PMDA approved drug
35807217|T121|Radiotherapy medication
35807218|T121|Topical
35807219|T121|Antiviral
35807220|T121|Irritant
35807221|T121|Antibody-drug conjugate
35807222|T121|Anti-HER2 antibody
35807223|T121|Microtubule inhibitor
35807224|T121|Mutation-specific medication
35807225|T121|EGFR inhibitor
35807226|T121|ERBB2 inhibitor
35807227|T121|ERBB4 inhibitor
35807228|T121|Cytokine
35807229|T121|ALK inhibitor
35807230|T121|Neutral
35807231|T121|Anti-CD52 antibody
35807232|T121|REMS program
35807233|T121|Bisphosphonate
35807187|T121|Aurora kinase inhibitor
35807234|T121|Retinoid
35807235|T121|WHO Essential Cancer Medicine
35807236|T121|Xanthine oxidase inhibitor
35807237|T121|Benzodiazepine
35807238|T121|Alkylating agent
35807239|T121|Orphan drug
35807240|T121|Anti-mesothelin antibody
35807241|T121|Chemotherapy protective agent
35807242|T121|Hematology medication
35807243|T121|Hemostasis medication
35807244|T121|Fibrinolysis inhibitor
35807245|T121|Aromatase inhibitor
35807246|T121|Intramuscular
35807247|T121|Antimetabolite
35807248|T121|Antifolate
35807249|T121|Discontinued drug
35807250|T121|Vesicant
35807251|T121|Human DNA synthesis inhibitor
35807252|T121|Health Canada approved drug
35807253|T121|Phosphodiesterase inhibitor
35807254|T121|Fractionated plasma product
35807255|T121|Coagulation factor
35807256|T121|Nonsteroidal antiandrogen
35807257|T121|VEGFR inhibitor
35807258|T121|KIT inhibitor
35807259|T121|SRC inhibitor
35807261|T121|Direct oral anticoagulant
35807262|T121|Factor Xa inhibitor
35807263|T121|Neurokinin 1 (NK1) antagonist
35807264|T121|Anticoagulant
35807265|T121|Direct thrombin inhibitor
35807266|T121|Subcutaneous
35807267|T121|Enzyme
35807268|T121|COX-1 inhibitor
35807269|T121|PDE inhibitor
35807270|T121|Anti-PD-L1 antibody
35807271|T121|Supportive medication
35807272|T121|Hematopoietic growth factor
35807273|T121|Megakaryocyte growth factor
35807274|T121|Cellular therapy
35807275|T121|PDGFR inhibitor
35807276|T121|Inflammitant
35807277|T121|Hypomethylating agent
35807278|T121|DNA methyltransferase inhibitor
35807279|T121|Pyrimidine analogue
35101588|T121|Chlorambusil
35101587|T121|Chloraminophene
35101586|T121|Chlorbutin
35807280|T121|Anti-DKK1 antibody
35101585|T121|Chlorobutin
35807281|T121|Immunotoxin
35807282|T121|Anti-CD22 antibody
35807283|T121|Halted drug
35807284|T121|Intravesical
35807285|T121|Anti-PS antibody
35807286|T121|Tumor vaccine
35807287|T121|KFDA approved drug
35807288|T121|Nitrogen mustard
35807289|T121|Anti-VEGFR antibody
35807290|T121|Biosimilar
35807291|T121|MAP2K1 inhibitor
35807292|T121|MAP2K2 inhibitor
35807293|T121|Intracavitary
35807294|T121|Anti-CD19 antibody
35807295|T121|Proteasome inhibitor
35807296|T121|Light-chain (AL) amyloidosis medication
35807297|T121|Bcr-Abl inhibitor
35807298|T121|Radiation
35807299|T121|Anti-CD30 antibody
35807300|T121|ROS1 inhibitor
35807301|T121|IGFR inhibitor
35807302|T121|FLT3 inhibitor
35807303|T121|PI3K inhibitor
35101584|T121|Chromo-Z
35807304|T121|Taxane
35807305|T121|AXL inhibitor
35807306|T121|MET inhibitor
35807307|T121|RET inhibitor
35807308|T121|TEK inhibitor
35807309|T121|TRK inhibitor
35807310|T121|Pegylated medication
35807311|T121|Mucositis prevention
35807312|T121|P2Y12 ADP inhibitor
35807313|T121|Fluoropyrimidine
35807314|T121|Anti-vWF medication
35807315|T121|Platinum agent
35807316|T121|Cancer of unknown primary medication
35807317|T121|Nitrosourea
35807318|T121|Intralesional
35807319|T121|Antifungal
35101583|T121|Cicoxil
35101582|T121|Cidaprim
35807320|T121|Anti-EpCAM antibody
35807321|T121|EMA approved drug
35807322|T121|Anti-PD-1 antibody
35807323|T121|Antihistamine
35807324|T121|Anti-EGFR antibody
35807325|T121|H2-receptor antagonist
35101581|T121|Cipaprim
35101580|T121|Ciplin
35101579|T121|Circuvit
35101578|T121|Citofolin
35101577|T121|Citosin
35101576|T121|Citrim
35101575|T121|Cladon
35807326|T121|Anti-IGF-1R antibody
35807327|T121|Purine analogue
35807328|T121|Antibacterial
35807329|T121|PI3K alpha inhibitor
35807330|T121|PI3K delta inhibitor
35807331|T121|Steroid
35807332|T121|Anti-P-selectin antibody
35807333|T121|Clusterin inhibitor
35807334|T121|Nasal
35807335|T121|Immunosuppressant
35101574|T121|Claro
35807336|T121|ciclosporin
35807336|T121|CsA
35807336|T121|cyclosporin
35807336|T121|cyclosporin A
35807336|T121|CyA
35807336|T121|Cyclosporine
35807337|T121|Calcineurin inhibitor
35807338|T121|Intrathecal
35101573|T121|Cleveron
35807339|T121|Deoxycytidine analogue
35807340|T121|Liposomal chemotherapy
35101572|T121|Clinitran
35101571|T121|Clonea
35807341|T121|BRAF inhibitor
35101570|T121|Clotrizol
35807342|T121|Triazene
35101569|T121|CO-Sultrin
35101568|T121|CO-Tasian
35101567|T121|CO-Traisole 480
35807343|T121|Heparin
35807344|T121|Low molecular weight heparin
35101566|T121|CO-Trim-Tablinen
35101565|T121|CO-Trimazole
35807345|T121|Anti-CD38 antibody
35101564|T121|CO-Trimed
35101563|T121|CO-Trimoxa
35101562|T121|CO-Trimoxazol
35807346|T121|Erythrocyte growth factor
35101561|T121|Cobact
35101560|T121|Cobal ST
35807347|T121|SYK inhibitor
35807348|T121|Chelator
35807349|T121|GnRH antagonist
35807350|T121|Anti-RANKL antibody
35807351|T121|RANK ligand inhibitor
35101559|T121|Cocydal
35807352|T121|Vasopressin analog
35101558|T121|Cofatrim
35807353|T121|Anti-GD2 antibody
35807354|T121|Laxative
35807355|T121|Serotonin 5-HT3 antagonist
35807356|T121|Dopamine receptor antagonist
35807357|T121|Phenothiazine
35807358|T121|FGFR inhibitor
35802853|T121|Intra-arterial
35807359|T121|Cannabinoid
35807360|T121|5 alpha-reductase inhibitor
35807361|T121|PI3K gamma inhibitor
35807362|T121|Anti-C5 antibody
35807363|T121|Anti-SLAMF7 antibody
35807364|T121|Bispecific antibody medication
35807365|T121|Anti-Factor IXa antibody
35807366|T121|Anti-Factor Xa antibody
35807367|T121|IDH2 inhibitor
35807368|T121|Adrenergic receptor agonist
35807369|T121|MTOR inhibitor
35807370|T121|TSC1 inhibitor
35807371|T121|TSC2 inhibitor
35807372|T121|Iron
35807373|T121|KSP inhibitor
35807374|T121|Granulocyte colony-stimulating factor
35807375|T121|WHO Essential Anti-infective Medicine
35807376|T121|Anabolic steroid
35807377|T121|Purine nucleoside phosphorylase (PNP) inhibitor
35807378|T121|Drugs PMDA approved in 2017
35807379|T121|Estrogen receptor inhibitor
35807380|T121|Diuretic
35807381|T121|Steroidal androgen receptor inhibitor
35807382|T121|Hsp90 inhibitor
35101557|T121|Colircusi Dexametasona
35101556|T121|Colitran
35807383|T121|Enediyne antibiotic
35101555|T121|Colizole
35807384|T121|Hedgehog pathway inhibitor
35807385|T121|GnRH agonist
35807386|T121|Antipsychotic
35807387|T121|Anti-CD47 antibody
35807388|T121|Anti-KIR antibody
35807389|T121|Anti-CD20 antibody
35807390|T121|Anti-CD20 medication
35807391|T121|Radioimmunoconjugate
35807392|T121|ITK inhibitor
35807393|T121|TEC inhibitor
35807394|T121|TXK inhibitor
35101554|T121|Colotrim
35807395|T121|Telomerase inhibitor
35807396|T121|COX-2 inhibitor
35807397|T121|Interferon
35807398|T121|Anti-CTLA-4 antibody
35101553|T121|Comax
35807399|T121|IDH1 inhibitor
35101552|T121|Comazole
35101551|T121|Combact
35807400|T121|Somatostatin analog
35807401|T121|Proton pump inhibitor
35101550|T121|Combi-Methoxan
35807402|T121|Anti-HER2 medication
35807403|T121|Immunomodulatory drugs (IMiDs)
35101549|T121|Comixco
35807404|T121|JAK inhibitor
35101548|T121|Comox
35807405|T121|Anti-diarrheal
35101547|T121|Comoxol
35807406|T121|Anti-TRAIL-R1 antibody
35807407|T121|PTK2 inhibitor
35807408|T121|Appetite stimulant
35807409|T121|Anti-IL-5 antibody
35807410|T121|Anti-CCR4 antibody
35807411|T121|Anti-CD194 antibody
35807412|T121|Antileukotriene
35807413|T121|Anti-amyloid antibody
35807414|T121|ERBB3 inhibitor
35807415|T121|ERBB2 (HER2) medication
35807416|T121|ERBB3 (HER3) medication
35807417|T121|CSF1R inhibitor
35807418|T121|DDR inhibitor
35807419|T121|PARP inhibitor
35807420|T121|Device
35807421|T121|Anti-PDGFR antibody
35807422|T121|Cephalotaxine
35807423|T121|Anti-c-Met antibody
35807424|T121|Anti-CD37 antibody
35807425|T121|Nanoparticle albumin bound chemotherapy
35101546|T121|Contrimoxazole
35807426|T121|MSI-H or dMMR medication
35807427|T121|Inhalation
35807428|T121|MEK inhibitor
35807429|T121|Drugs EMA approved in 2013
35807430|T121|CXCR4 inhibitor
35807431|T121|Alpha emitter
35807432|T121|Selective estrogen receptor modulator
35807433|T121|Uric acid lowering agent
35807434|T121|Anti-HGF antibody
35807435|T121|Anti-TACSTD2 antibody
35807436|T121|Granulocyte macrophage colony-stimulating factor
35807437|T121|Muscarinic receptor antagonist
35807438|T121|XPO1 inhibitor
35807439|T121|Ultralow molecular weight heparin
35807440|T121|Anti-IL-6 antibody
35807441|T121|Dendritic cell vaccine
35807442|T121|SMO inhibitor
35807443|T121|Intervention index
35807444|T121|Oncolytic viral therapy
35807445|T121|Tryptophan hydroxylase inhibitor
35807446|T121|Anti-TRAIL-R2 antibody
35807447|T121|Farnesyltransferase inhibitor
35807448|T121|Chimeric antigen receptor T-cell
35101545|T121|Coprim
35101544|T121|Coprime
35807449|T121|Anti-IL-6R antibody
35807450|T121|Aminopeptidase inhibitor
35807451|T121|Peptibody medication
35807452|T121|Anti-CD27 antibody
35807453|T121|MAP2K4 inhibitor
35807454|T121|MAP3K20 inhibitor
35807455|T121|MAP4K5 inhibitor
35807456|T121|Bcl-2 inhibitor
35807457|T121|Vinca alkaloid
35807460|T121|SMO or PTCH-1 (Hedgehog) medication
35807461|T121|PLK1 inhibitor
35807462|T121|PAR1 inhibitor
35807463|T121|Vitamin K antagonist
35807464|T121|Soluble decoy receptor
42542303|T121|Autoimmune hematologic condition
42542304|T121|Bleeding disorder
42542305|T121|Acute leukemia
42542306|T121|Endocrine cancer
35101543|T121|Corodex
42542307|T121|T-cell lymphoma
42542308|T121|Gastrointestinal cancer
42542309|T121|High-grade glioma
42542310|T121|Thrombotic disorder
42542311|T121|Bone marrow failure syndrome
42542312|T121|Cytopenia
42542313|T121|Complementopathy
42542314|T121|Pediatric cancer
42542315|T121|Genitourinary cancer
42542316|T121|Aggressive lymphoma
42542317|T121|Non-Hodgkin lymphoma
42542318|T121|CNS cancer
42542319|T121|Lymphoproliferative disorder
42542320|T121|Gynecologic cancer
42542321|T121|Hepatobiliary cancer
42542322|T121|Indolent lymphoma
42542323|T121|Myeloproliferative neoplasm
42542324|T121|Colorectal cancer
42542325|T121|Cutaneous lymphoma
42542326|T121|Non-melanoma skin cancer
42542327|T121|Histiocytosis
42542328|T121|Alloimmune hematologic condition
42542329|T121|Plasma cell dyscrasia
42542330|T121|Skin cancer
42542331|T121|Thoracic cancer
42542332|T121|Lung cancer
42542333|T121|Inherited hemoglobinopathy
42542334|T121|T-cell leukemia
35802854|T121|Drug
35807465|T121|Intervention
35807466|T121|Antineoplastics by class effect
35807467|T121|Routed medication
35807468|T121|Antiplatelet agent
35807469|T121|Biomarker-specific medication
35807470|T121|Site-specific medication
35807471|T121|Enzyme inhibitor
35807472|T121|Malignant hematology medication
35807473|T121|Genitourinary oncology medication
35807474|T121|Approved drug
35807475|T121|WHO Essential Medicine
35807476|T121|Antibiotic
35807477|T121|Thoracic oncology medication
35807478|T121|Growth factor inhibitor
35101542|T121|Corson
35101541|T121|Corsona
35101540|T121|Corsone
35101539|T121|Corsum
35807479|T121|Pediatric oncology medication
35807480|T121|Classical hematology medication
35807481|T121|Bone protective medication
35807482|T121|Gynecologic oncology medication
35807483|T121|Biologic product
35807484|T121|Coagulopathy medication
35807485|T121|Gastrointestinal oncology medication
35807486|T121|Thrombosis medication
35101538|T121|Cortesa
35807487|T121|Nonsteroidal anti-inflammatory drugs (NSAIDs)
35807488|T121|Endocrine oncology medication
35101537|T121|Corticoidex
35101536|T121|Cortidax
35101535|T121|Cortidex
35807489|T121|Site-agnostic medication
35101534|T121|Cortidexason
35807490|T121|Neurooncology medication
35101533|T121|Cortisolona
35101532|T121|Cortitop
35807491|T121|Drugs by vehicle
35807492|T121|Histiocytoses medication
35101531|T121|Cosat
35807493|T121|Immunosuppresant
35807494|T121|Molecular chaperone inhibitor
35807495|T121|Bowel management
35807496|T121|GTPase-activating protein inhibitor
35807497|T121|Granulocyte growth factor
35807498|T121|Drugs PMDA approved in the 2010'
35807499|T121|Drugs PMDA approved in the 21st century
35101530|T121|Cosig
35807500|T121|Androgen receptor inhibitor
35807501|T121|Drugs EMA approved in the 2010'
35807502|T121|Drugs EMA approved in the 21st century
35807503|T121|Selective inhibitors of nuclear export
35807504|T121|Immune effector cell
35807505|T121|Apoptosis promoter
42542335|T121|Classical hematologic condition
42542336|T121|Malignant hematologic neoplasm
42542337|T121|Lymphoma
42542338|T121|T-cell neoplasm
42542339|T121|Cross-disciplinary condition
42542340|T121|Hemoglobinopathy
42542341|T121|Leukemia
42542342|T121|Sarcoma
35807506|T121|Pre-definitive therapy
35807507|T121|Post-definitive therapy
35101529|T121|Costazole
35807508|T121|Curative therapy
35807509|T121|Non-curative second-line induction therapy
35101528|T121|Cosulf
35807510|T121|Non-curative third-line induction therapy
35807511|T121|Non-curative third-line consolidation therapy
35807512|T121|Non-curative third-line maintenance therapy
35807513|T121|Non-curative subsequent-line induction therapy
35101527|T121|ADT and Darolutamide
35101526|T121|Anti-diarrheals
35101525|T121|Anti-IFNg antibody
35101524|T121|Anticoagulants
35101523|T121|Antiplatelet agents
35101522|T121|Ascorbic acid
35101521|T121|Atarax
35101520|T121|Bendamustine and Brentuximab vedotin
35101520|T121|Brentuximab Vedotin and Bendamustine
35101519|T121|Bilateral salpingo-oophorectomy
35101518|T121|Clonazepam
35101517|T121|Cyclosporine and Mycophenolate mofetil
35101516|T121|Cyclosporine, Mycophenolate mofetil, Sirolimus
35101515|T121|NI-0501
35101515|T121|emapalumab-lzsg
35101515|T121|Emapalumab
35101514|T121|Gamifant
35101513|T121|Hydroxyzine
35101512|T121|Klonopin
35101511|T121|Meperidine
35101510|T121|Nonsteroidal androgen receptor inhibitors
35101509|T121|Nubeqa
35101508|T121|RBC transfusions
42542343|T121|Pentostatin and Alemtuzumab
42542344|T121|GemOx and Sorafenib
42542344|T121|Gemcitabine, Oxaliplatin , Sorafenib
42542345|T121|mFOLFOX and Sorafenib
42542345|T121|modified FOLinic acid, Fluorouracil, OXaliplatin, Sorafenib
42542346|T121|HAIC and Sorafenib
35101507|T121|AC-T
35101507|T121|Adriamycin (Doxorubicin) and Cyclophosphamide followed by Taxol (Paclitaxel)
35101506|T121|Acic
35101505|T121|Aciphex
35101504|T121|Acivir
35101503|T121|Acivirax
35101502|T121|Actemra
35101501|T121|Actimmune
35101500|T121|Actonel
35101499|T121|Acylete
35101498|T121|Amixam
35101497|T121|Ammoidin
35101496|T121|Amoxi
35101495|T121|Amoxihexal
35101494|T121|Amoxil
35101493|T121|Anastrozole and Palbociclib
35101492|T121|Andexxa
35101491|T121|Androcur
35101490|T121|Apo-acyclovir
35101489|T121|Avorax
35101488|T121|Axcel
35101487|T121|Binorel
35101486|T121|Biomox
35101485|T121|Biovelbin
35101484|T121|Brilinta
35101483|T121|Brilique
35101482|T121|CALGB 8811 early intensification
35101481|T121|CALGB 8811 late intensification
35101990|T121|Capecitabine and Fulvestrant
35101989|T121|Caphosol
35101988|T121|CHVmP
35101987|T121|CHVmP-VB
35101987|T121|Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Vm26 (Teniposide), Prednisone, Vincristine, Bleomycin
35101986|T121|Cyclophosphamide and Methotrexate (CM)
35101986|T121|CM
35101986|T121|Cyclophosphamide and Methotrexate
42542347|T121|AV-CMF
42542348|T121|AVCF
42542348|T121|Adriamycin (Doxorubicin), Vincristine, Cyclophosphamide, Fluorouracil
42542349|T121|Calaspargase, Daunorubicin, Vincristine, Prednisone
42542350|T121|Carboplatin and Cyclophosphamide
42542351|T121|CAV and RT
42542351|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Vincristine, Radiation Therapy
42542352|T121|CAVE
42542352|T121|CAV-E
42542352|T121|Cyclophosphamide, Adriamycin (Doxorubicin), Vincristine, Etoposide
42542353|T121|CEV (Cyclophosphamide/Etoposide)
42542353|T121|CEV
42542353|T121|Cyclophosphamide, Etoposide, Vincristine
42542354|T121|Dose-dense Epirubicin monotherapy
42542354|T121|dose-dense Epirubicin
42542355|T121|Docetaxel and Nintedanib
42542356|T121|EMA-CO
42542356|T121|Etoposide, Methotrexate, Actinomycin D, Cyclophosphamide, Oncovin (Vincristine)
42542357|T121|Etoposide, Ifosfamide, Imatinib
42542358|T121|Euflex
42542359|T121|FCR (Rituximab and hyaluronidase)
42542359|T121|Fludarabine, Cyclophosphamide, Rituximab hyaluronidase
42542360|T121|FUIRI
42542360|T121|5-FU and IRInotecan
42542361|T121|FULV and Bevacizumab
42542361|T121|5-FU, LeucoVorin (Folinic acid), Bevacizumab
42542362|T121|FUOX
42542362|T121|5-FU and OXaliplatin
42542363|T121|Histrelin monotherapy
42542364|T121|Hydroxyurea and Plicamycin
42542365|T121|Cyclophosphamide, Mycophenolate mofetil, Tacrolimus
42542366|T121|Lomustine and Bevacizumab
42542367|T121|Methotrexate and Tacrolimus
42542368|T121|Mitoxantrone and Hydrocortisone
42542369|T121|Nintedanib and Pemetrexed
42542370|T121|Ofev
42542371|T121|Pegaspargase, Vincristine, Prednisone
42542372|T121|PUVA
42542372|T121|Psoralen and Ultra-Violet A
42542373|T121|R-CHOP-14 (Rituximab and hyaluronidase)
42542373|T121|Rituximab and hyaluronidaase, Cyclophosphamide, Hydroxydaunorubicin (Doxorubicin), Oncovin (Vincristine), Prednisone every 14 days
42542374|T121|Rituximab and hyaluronidase monotherapy
42542375|T121|STAMP-I
42542376|T121|Carboplatin and Paclitaxel (CP) and Nintedanib
42542376|T121|CP and Nintedanib
42542376|T121|TC and Nintedanib
42542376|T121|Carboplatin, Paclitaxel, Nintedanib
42542376|T121|Taxol (Paclitaxel), Carboplatin, Nintedanib
42542377|T121|VAB-6
42542378|T121|Valrubicin monotherapy
42542379|T121|Vargatef
42542380|T121|IVIG monotherapy
42542381|T121|Kanjinti
42542382|T121|Lenvatinib and Pembrolizumab
42542383|T121|Ontruzant
42542384|T121|Prednisolone and Rituximab
42542385|T121|Prednisone and Rituximab
42542386|T121|Rituximab-pvvr
42542387|T121|Ruxience
42542388|T121|Trastuzumab-anns
42542389|T121|Trastuzumab-dttb
42542390|T121|Trastuzumab-qyyp
42542391|T121|Trazimera
35101985|T121|Cusiviral
35101984|T121|Cyclophosphamide, Cytarabine, Pegaspargase, Thioguanine, Vincristine, Dexamethasone
35101983|T121|Cyclovax
35101982|T121|Cyclovir
35101981|T121|Cyklokapron
35101980|T121|Cytomega
35101979|T121|Dara-KD
35101978|T121|Dose-dense AC-T
35101978|T121|ddAC-T
35101978|T121|dose-dense Adriamycin (Doxorubicin) and Cyclophosphamide followed by Taxol (Paclitaxel)
35101977|T121|Declovir
35101976|T121|Deltasoralen
35101975|T121|Demerol
35101974|T121|Depacon
35101973|T121|Depakine
35101972|T121|Depakote
35101971|T121|Dermox
35101970|T121|Desplex
35101969|T121|Dibestrol
35101968|T121|Dilantin
35101967|T121|Dravyr
35101966|T121|Ductaclose
35101965|T121|Elmetacin
35101964|T121|Encorate
35101963|T121|Entrectinib monotherapy
35101962|T121|Epanutin
35101961|T121|Epibest
35101960|T121|Epilim
35101959|T121|Epival
35101958|T121|Epsotoin
35101957|T121|Eptoin
35101956|T121|Eunades
912154|T121|Everolimus and Vinorelbine
35101955|T121|Evista
35101954|T121|Ex-Lax
35101953|T121|SAR302503
35101953|T121|TG101348
35101953|T121|Fedratinib
35101952|T121|Fedratinib monotherapy
35101951|T121|Fentinol
35101950|T121|Flonorbin
35101949|T121|Gemcitabine and Trastuzumab
35101948|T121|Geralen
35101947|T121|Geroxalen
35101946|T121|Hemostan
35101945|T121|Hepirax
35101944|T121|Herceptin Hylecta
35101943|T121|Herpevex
35101942|T121|Herpex
35101941|T121|Herzovir
35101940|T121|Hycamtin
35101939|T121|Indocid
35101938|T121|Indocin
35101937|T121|Indocrom
35101936|T121|Indoga
35101935|T121|Inmecin
35101934|T121|Inrebic
35101933|T121|Irinotecan and S-1
35101932|T121|Javlor
35101931|T121|Klovireks-l
35101930|T121|Leeporate
35101480|T121|Lentaron
35101479|T121|Lovir
35101478|T121|Lucanix
35101477|T121|LymphoCide
35101476|T121|Medovir
35101475|T121|Meladinina
35101474|T121|Meladinine
35101473|T121|Mercaptopurine, Methotrexate, Vincristine, Dexamethasone
35101472|T121|Metastron
35101471|T121|Methotrexate and Pegaspargase
35101470|T121|Metoxaleno
35101469|T121|Mithracin
35101468|T121|Mopsoralen
35101467|T121|nab-Paclitaxel and Trastuzumab
35101466|T121|Navelbine
35101465|T121|Neoben
35101464|T121|Neumega
35101463|T121|Nidran
35101462|T121|Nilevar
35101461|T121|Nplate
35101460|T121|Nublexa
35101459|T121|Ogivri
35101457|T121|Orafix
35101456|T121|Ortrex
35101455|T121|Orvor
35101454|T121|Oxsoralen
35101453|T121|Oxsoralen-Ultra
35101452|T121|Paclitaxel and Vinorelbine
35101451|T121|Paclitaxel, Pertuzumab, Ado-trastuzumab emtansine
35101451|T121|Paclitaxel, Pertuzumab, Trastuzumab emtansine
35101286|T121|Pariet
35101285|T121|Perdiem
35101284|T121|Pharmaniaga
35101458|T121|Photofrin
35101283|T121|Prexam
35101282|T121|Puvasoralen
35101281|T121|Qualaquin
35101280|T121|Quizartinib monotherapy
35101279|T121|Rablet
35101278|T121|Ralista
35101277|T121|Razylan
35101276|T121|Reconaz
35101275|T121|Regonix
35101274|T121|Relbovin
35101273|T121|Removab
35101272|T121|Renib
35101271|T121|Resihance
35101270|T121|RhoGAM
35101269|T121|Ribone
35101268|T121|Risedol
35101267|T121|Risofos
35101266|T121|Rituxan Hycela
35101265|T121|Rozlytrek
35101264|T121|Saforax
35101263|T121|Senokot
35101262|T121|SOX and Bevacizumab
35101262|T121|S-1, OXaliplatin, Bevacizumab
35101261|T121|Stibrol
35101260|T121|Stilbest
35101259|T121|Stivarga
912155|T121|TEC
35101258|T121|Temsy
35101257|T121|Ticalog
35101256|T121|Tivorbex
35101255|T121|Topecan
35101254|T121|Topotec
35101253|T121|Tranofast
35101252|T121|trastuzumab and hyaluronidase-oysk
35101252|T121|Trastuzumab and hyaluronidase
35101251|T121|Ultramop
35101250|T121|Uvadex
35101249|T121|V-Gavir
35101248|T121|Vacrax
35101247|T121|VagaCyte
35101246|T121|Valcyclovir
35101245|T121|Valcyte
35101244|T121|Valgan
35101243|T121|Valixa
35101242|T121|Vallona
35101241|T121|Valnov
35101240|T121|Valric
35101239|T121|Valstar
35101238|T121|Valtaxin
35101237|T121|Verz
35101236|T121|Vfend
35101235|T121|Vicide
35101234|T121|Vinelbine
35101233|T121|Vinorelbel
35101232|T121|Vinotec
35101231|T121|Virax
35101230|T121|Virest
35101229|T121|Virless
35101228|T121|Virolfi
35101227|T121|Virox
35101226|T121|Virucid
35101225|T121|Virupos
35101224|T121|Vonaz
35101223|T121|Voraze
35101222|T121|Voricort
35101221|T121|Vorier
35101220|T121|Vorirx
35101219|T121|Voritek
35101218|T121|Voritrol
35101217|T121|Voriva
35101216|T121|Vorizol
35101215|T121|Vorwell
35101214|T121|Vorzole
35101213|T121|Vorzu
35101212|T121|Welldom
35101211|T121|Xanthotoxin
35101210|T121|Xovir
35101209|T121|Zantac
35101208|T121|Zarnestra
35101207|T121|Zevin
35101206|T121|Zirax
35101205|T121|Zoral
35101204|T121|Zorax
35101203|T121|Zoraxin
35101202|T121|Zoviax
35101201|T121|Zovir
35101200|T121|Zovirax
42542392|T121|Melphalan, then Fludarabine, Busulfan, ATG, then allo HSCT
42542393|T121|Anakinra monotherapy
42542394|T121|Binimetinib, Encorafenib, Cetuximab
42542395|T121|BRAF-mutated Colorectal cancer
42542396|T121|Carboplatin and Etoposide (CE) and Durvalumab
42542397|T121|CCI
42542397|T121|Cisplatin, Carboplatin, Ifosfamide
42542398|T121|Cisplatin and Etoposide (EP) and Durvalumab
42542399|T121|Cisplatin, Fluorouracil, Pembrolizumab
42542400|T121|Cisplatin, Pemetrexed, TTFields
42542401|T121|Colchicine monotherapy
42542402|T121|Crizanlizumab monotherapy
42542403|T121|Dabrafenib, Trametinib, Panitumumab
912156|T121|EP and Ipilimumab
912157|T121|EP, Tamoxifen, RT
42542404|T121|Erlotinib and Ramucirumab
42542405|T121|Interferon alfa-n1 monotherapy
42542406|T121|Irinotecan, Vemurafenib, Cetuximab
42542407|T121|Pomalidomide and Dexamethasone (PD)
42542407|T121|Pomalidomide and low-dose dexamethasone
912158|T121|PD and Pembrolizumab
42542408|T121|Pipobroman monotherapy
42542409|T121|T-cell prolymphocytic leukemia
42542410|T121|TILs
42542410|T121|Tumor Ifiltrating Lymphocytes
42542411|T121|BGB-3111
42542411|T121|Zanubrutinib
42542412|T121|Zanubrutinib monotherapy
42542413|T121|Anthracycline-containing regimen
42542414|T121|Bevacizumab-containing regimen
42542415|T121|Irinotecan-containing regimen
42542416|T121|IRIS
42542417|T121|Platinum doublet
42542418|T121|Anti-Factor XIa antibody
42542419|T121|Antiestrogen-containing regimen
42542420|T121|ABL001
42542420|T121|Asciminib
42542421|T121|BRCA-mutated Ovarian cancer
42542422|T121|BRCA-mutated Pancreatic cancer
42542423|T121|Epithelioid sarcoma
42542424|T121|Erythropoietin monotherapy
42542425|T121|EZH2 inhibitor
42542426|T121|Fluorouracil and Paclitaxel
42542427|T121|Giant-cell tumor of bone
42542428|T121|HER2-positive - historical Breast cancer
42542429|T121|HER2-positive Colorectal cancer
42542430|T121|Intron-A
42542431|T121|Kaposi sarcoma
42542432|T121|KIT-mutated Melanoma
42542433|T121|KRAS-mutated Non-small cell lung cancer
42542434|T121|Leiomyosarcoma
42542435|T121|Liposarcoma
42542436|T121|ACE-536
42542436|T121|luspatercept-aamt
42542436|T121|Luspatercept
42542437|T121|Luspatercept monotherapy
42542438|T121|BAY 1213790
42542438|T121|Osocimab
42542439|T121|Reblozyl
42542440|T121|Rituximab-containing regimen
42542441|T121|E7438
42542441|T121|EPZ6438
42542441|T121|Tazemetostat
42542442|T121|Tazemetostat monotherapy
42542443|T121|Tazverik
42542444|T121|TCHP (Paclitaxel)
42542444|T121|TCHP
42542444|T121|Taxol (Paclitaxel), Carboplatin, Herceptin (Trastuzumab), Pertuzumab
42542445|T121|Teniposide and WBRT
42542446|T121|Triptorelin monotherapy
42542447|T121|Vepesid
912159|T121|ICE and ATRA
912159|T121|Idarubicin, Cytarabine, Etoposide, All-Trans Retinoic Acid
912160|T121|Immunostimulatory monoclonal antibody
912161|T121|Immunosuppressive monoclonal antibody
912162|T121|NPM1-mutated Acute myeloid leukemia
912163|T121|Targeted therapeutic
912164|T121|Viral DNA synthesis inhibitor
912165|T121|Imuran
912166|T121|Indenza
912167|T121|Interferon alfa-2c
912168|T121|Interferon alfa-n1
912169|T121|KRAS inhibitor
912170|T121|KRD-PACE
912170|T121|Kyprolis (Carfilzomib), Revlimid (Lenalidomide), Dexamethasone, Platinol (Cisplatin), Adriamycin (Doxorubicin), Cyclophosphamide, Etoposide
912171|T121|Kryxana
912174|T121|Litican
912175|T121|Lucicaboz
912176|T121|Lucicer
912177|T121|Lucipalb
912178|T121|Margenza
912179|T121|MGAH22
912179|T121|Margetuximab
912180|T121|Mitigare
912181|T121|Mostarina
912172|T121|Noxalk
912173|T121|Ocular adenexal MALT lymphoma, antibiotic therapy
912182|T121|Orgovyx
912183|T121|Palbace
912184|T121|Palbocap
912185|T121|Palbocent
912186|T121|Palbonix
912187|T121|Plenaxis
912188|T121|Quinamed
912189|T121|RAF1 inhibitor
912190|T121|Relumina
912191|T121|Serine-threonine kinase inhibitor
912192|T121|Sitagliptin, Sirolimus, Tacrolimus
912193|T121|AMG 510
912193|T121|Sotorasib
912194|T121|Spexib
912195|T121|Sterocyt
912196|T121|Tauritmo
912197|T121|Trepmac
912198|T121|Tyrosine kinase inhibitor
912199|T121|TGR-1202
912199|T121|Umbralisib
912200|T121|Vercite
912201|T121|Vercyte
912202|T121|Verzenios
912203|T121|WEE1 inhibitor
912204|T121|Xanafide
35101199|T121|Cotoram
912205|T121|ME
35101198|T121|Cotran
35101197|T121|Cotrazen
912206|T121|AME
912207|T121|A-ICE
912208|T121|FLAI
35101196|T121|Cotrexel
912209|T121|FLA
912210|T121|VADx
35101195|T121|Cotri
912211|T121|Cytarabine and Vosaroxin
35101194|T121|Cotribase
35101193|T121|Cotribene
35101192|T121|Cotribid
35101191|T121|Cotril
35101190|T121|Cotrilin
912212|T121|CAD
35101189|T121|Cotrim
912213|T121|FAP
35101188|T121|Cotrimax
35101187|T121|Cotrimaxazol
912214|T121|Epirubicin and Vinorelbine (VE)
912214|T121|VE
912214|T121|Vinorelbine and Epirubicin
35101186|T121|Cotrimaxazole
35807514|T121|Oopherectomy
35101185|T121|Cotrimel
35101184|T121|Cotrimhexal
35101183|T121|Cotrimol
35101182|T121|Cotrimox
35101181|T121|Cotrimoxazol
35101180|T121|Cotrimoxin
35101179|T121|Cotrimstada
35101178|T121|Cotripharm
35101177|T121|Cotrisul
35807515|T121|Surgery
35101176|T121|Cotrixyl-L
912215|T121|AC-TL (Paclitaxel)
912215|T121|AC-TL
912215|T121|"<div class=""toccolours"" style=""background-color:#eeeeee"">"
912215|T121|Adriamycin (Doxorubicin) and Cyclophosphamide, followed by Taxol (Paclitaxel) and Lapatinib
35101175|T121|Cotrizol
912216|T121|MTP
35101174|T121|Cotrizole
912217|T121|Afatinib and Vinorelbine
35101173|T121|Cots
912218|T121|3M
912219|T121|VNC
912220|T121|CIB
912221|T121|MMF
912222|T121|MFL
912223|T121|FOLF-CB
912224|T121|ECVBP
35101172|T121|Coumadin
35101171|T121|Coumadine
35807516|T121|Surgery alone
912225|T121|PELF
912226|T121|EAP
35101170|T121|Couparin
912227|T121|FA
912227|T121|Fluorouracil and Adriamycin (Doxorubicin)
912228|T121|ELF
912229|T121|VAPEC-B
911922|T121|TPCV
912230|T121|VCE
912231|T121|VBD
912232|T121|DBCT
912233|T121|VTDC
912234|T121|Bortezomib and Bevacizumab
912235|T121|Bortezomib and Siltuximab
912236|T121|MPP
912237|T121|Carboplatin and Paclitaxel (CP) and Erlotinib
912238|T121|Carboplatin and Paclitaxel (CP) and Bexarotene
912239|T121|Carboplatin and Paclitaxel (CP) and Sorafenib
912240|T121|Carboplatin and Paclitaxel (CP) and Cediranib
912241|T121|CP and Veliparib
912242|T121|CP and Cetuximab
912243|T121|NIP
912244|T121|Pemetrexed and Vandetanib
912245|T121|Pemetrexed and Cetuximab
912246|T121|CCG
912247|T121|CarboMIP
912248|T121|MEV
912249|T121|MVC
912250|T121|TCG
912251|T121|Carboplatin and Epirubicin
912252|T121|Carboplatin and Topotecan
912253|T121|Cisplatin and Gemcitabine (GC) and Cetuximab
35807517|T121|Bilateral orchiectomy
912254|T121|Vinorelbine and Hydrocortisone
35807518|T121|Deferred orchiectomy
912255|T121|Carboplatin and Etoposide (CE) and Ipilimumab
912256|T121|PEI
912257|T121|BTOC
912258|T121|CODE
912259|T121|CYVADIC
912260|T121|VPV
912261|T121|BV
35807519|T121|Null therapy
35807520|T121|Antibiotic therapy
35807521|T121|Tumor treating fields
35807522|T121|Antifibrinolytic therapy
35101169|T121|Coyensu
35101168|T121|Cozol
35101167|T121|Cozole
35101166|T121|Creptrim
35101165|T121|Cromatonbic Folinico
35101164|T121|Curaprim
35101163|T121|Cysplatyna
35101162|T121|Cytoferon
35101161|T121|D-Cort
35101160|T121|Dacrosone
35101159|T121|Dagonal
35101158|T121|Daidoron
35101157|T121|Daiphen
35101156|T121|Dalalone
35101155|T121|Dalisol
35101154|T121|Danason
35101153|T121|Danasone
35101152|T121|Danofran
35101151|T121|Dantenk
35101150|T121|Dara-VTD
35101150|T121|D-VTD
35101150|T121|Daratumumab, Velcade (Bortezomib), Thalidomide, Dexamethasone
35101149|T121|Daxilone
35101148|T121|Deca Forte
35101147|T121|Decacin
35101146|T121|Decacort
35101145|T121|Decaderm
35101144|T121|Decadolone
35101143|T121|Decadran
35101142|T121|Decadron
35101141|T121|Decadronal
35101140|T121|Decadronfosfat
35101139|T121|Decafos
35101138|T121|Decalin
35101137|T121|Decalon
35101136|T121|Decalona
35101135|T121|Decan
35101134|T121|Decans
35101133|T121|Decaron
35101132|T121|Decason
35101131|T121|Decasone
35101130|T121|Decaspray
35101129|T121|Decatrim
35101128|T121|Decazol
35101127|T121|Decdak
35101126|T121|Decdan
35101125|T121|Decicort
35101124|T121|Decilone
35101123|T121|Decobel
35101122|T121|Decolite
35101121|T121|Decone
35101120|T121|Decordex
35101119|T121|Decorex
35101118|T121|Decoron
35101117|T121|Decorten
35101116|T121|Dectan
35101115|T121|Dectancyl
35101114|T121|Deexa
35101113|T121|Defibrotide monotherapy
35101112|T121|Defixal
35101111|T121|Deflaren
35101110|T121|Degalin
35101109|T121|Dekesu
35101108|T121|Dekisachosei
35101107|T121|Dekort
35101106|T121|Deksa
35101105|T121|Deksalon
35101104|T121|Deksamet
35101103|T121|Dellamethasone
35101102|T121|Deltafluorene
35101101|T121|Demasone
35101713|T121|Demeson
35101712|T121|Denfos
35101711|T121|Deotrim
35101710|T121|Depmedalone
35101709|T121|Depo Melcort
35101708|T121|Depo Moderin
35101707|T121|Depo-Medrate
35101706|T121|Depo-Medrol
35101705|T121|Depoject
35101704|T121|Depomedrone
35101703|T121|Deposet
35101702|T121|Dermadex
35101701|T121|Dermidron
35101700|T121|Deron S
35101699|T121|Deronil
35101698|T121|Derson
35101697|T121|Dersone
35101696|T121|Dertrin
35101695|T121|Desalark
35101694|T121|Desametasone Fosf
35101693|T121|Desason
35101692|T121|Deson
35101691|T121|Detametazon
35101690|T121|Detasone
35101689|T121|Dethamedin
35101688|T121|Dexa
35101687|T121|Dexa Clinit
35101686|T121|Dexabene
35101685|T121|Dexabeta
35101684|T121|Dexacen-4
35101683|T121|Dexacilin
35101682|T121|Dexacip
35101681|T121|Dexacollyre
35101680|T121|Dexacom
35101679|T121|Dexacort
35101678|T121|Dexacortal
35101677|T121|Dexacortin
35101676|T121|Dexacortisone
35101675|T121|Dexacortisyl
35101674|T121|Dexacotsil
35101673|T121|Dexacron
35101672|T121|Dexacutis
35101671|T121|Dexaden
35101670|T121|Dexaderm
35101669|T121|Dexaderme
35101668|T121|Dexadermil
35101667|T121|Dexadon
35101100|T121|Dexadrol
35101099|T121|Dexadron
35101098|T121|Dexaedo
35101097|T121|Dexafar
35101096|T121|Dexafarm
35101095|T121|Dexaflam
35101094|T121|Dexaflan
35101093|T121|Dexagalen
35101092|T121|Dexagee
35101091|T121|Dexagel
35101090|T121|Dexagenta
35101089|T121|Dexaglos
35101088|T121|Dexagreen
35101087|T121|Dexagrin
35101086|T121|Dexahexal
35101085|T121|Dexaleniens
35101084|T121|Dexalocal
35101083|T121|Dexaltin
35101082|T121|Dexamag
35101081|T121|Dexamark
35101080|T121|Dexame
35101079|T121|Dexamecortin
35101078|T121|Dexamedis
35101077|T121|Dexamedix
35101076|T121|Dexamedron
35101075|T121|Dexameral
35101074|T121|Dexameson
35101073|T121|Dexamesone
35101072|T121|Dexamet
35101071|T121|Dexametason
35100968|T121|Dexametasona
35100967|T121|Dexametax
35100966|T121|Dexametazon
35100965|T121|Dexametazona
35100964|T121|Dexameth
35100963|T121|Dexamethason
35100962|T121|Dexamethasonum
35100961|T121|Dexamethazon
35100960|T121|Dexamethazone
35100959|T121|Dexametin
35100958|T121|Dexametisona
35100957|T121|Dexametonal
35100956|T121|Dexametrat
35100955|T121|Dexamex
35100954|T121|Dexamil
35100953|T121|Dexamine
35100952|T121|Dexaminor
35100951|T121|Dexamo
35100950|T121|Dexamonozon N
35100949|T121|Dexan
35100948|T121|Dexanel
35100947|T121|Dexanil
35100946|T121|Dexano
35100945|T121|Dexaphos
35100944|T121|Dexapolcort
35100943|T121|Dexapro
35100942|T121|Dexaril
35100941|T121|Dexaroid
35100940|T121|Dexaron
35100939|T121|Dexart
35100938|T121|Dexasin
35100937|T121|Dexasine
35100936|T121|Dexasol
35100935|T121|Dexasolone
35100934|T121|Dexason
35100933|T121|Dexasone
35100932|T121|Dexasonlin
35100931|T121|Dexatab
35100930|T121|Dexaton
35100929|T121|Dexatop
35100928|T121|Dexatotal
35100927|T121|Dexaval
35100926|T121|Dexaven
35100925|T121|Dexavet
35100924|T121|Dexawal
35100923|T121|Dexawieb
35100922|T121|Dexazen
35100921|T121|Dexazona
35100920|T121|Dexazone
35100919|T121|Dexicorta
35100918|T121|Dexin
35100917|T121|Dexinga
35100916|T121|Dexion
35100915|T121|Dexmene
35100914|T121|Dexmesone
35100913|T121|Dexmetha
35100912|T121|Dexmethasone
35100911|T121|Dexmethsone
35100910|T121|Dexona
35100909|T121|Dexone
35100908|T121|Dexonium
35100907|T121|Dexoptic
35100906|T121|Dexpak
35100905|T121|Dexsol
35100904|T121|Dexstar
35100903|T121|Dextason
35100902|T121|Dexthasol
35100901|T121|Dexton
35100900|T121|Dextrasone
35100899|T121|Dhatrin
35100898|T121|Dicorsone
35100897|T121|Dicosheun
35100896|T121|Dino-BAC
35100895|T121|Diometa
35100894|T121|Diseptyl
35100893|T121|Dison
35100892|T121|Dispred
35100891|T121|Divifolin
35100890|T121|DM Solone
35100889|T121|Doctrim
35100888|T121|Donray
35100887|T121|Dorison
35100886|T121|Doronil
35100885|T121|Dosatran
35100884|T121|Doxorubicin, Mercaptopurine, Pegaspargase, Vincristine, Prednisolone
35100883|T121|Drate
35100882|T121|Drenex
35100881|T121|Drilozole
35100880|T121|Dronadil
35100879|T121|Dronal
35100878|T121|Dronalent
35100877|T121|Dronat
35100876|T121|Drossul
35100875|T121|Drovitan
35100874|T121|Droxol
35100873|T121|Drxaline
35100872|T121|Drylin
35100871|T121|Dubac
35100870|T121|Dumotrim
35100869|T121|DUO Septol
35100868|T121|Duobact
35100867|T121|Duobiocin
35100866|T121|Duoctrin
35100865|T121|Duralone
35100864|T121|Duratrimet
35100863|T121|Durofolin
35100862|T121|Durost
35100861|T121|Dutran
35100860|T121|Duvaxan
35100859|T121|Dvaseptol
35100858|T121|Dynaprim
35100857|T121|Ecofol
35100856|T121|Ectaprim
35100855|T121|Ectrin
35100854|T121|Editrim
35100853|T121|Eduprim
35100852|T121|Egiferon
35100851|T121|Elandur
35100850|T121|Eliprim
35100849|T121|Elixirmethasone
35100848|T121|Elvefocal
35100847|T121|Emeran
35100846|T121|Emeset
35100845|T121|Emetra
35100844|T121|Emetron
35100843|T121|Emigo
35100842|T121|Emistat
35100841|T121|Emivox
35100840|T121|Emovis
35100839|T121|Endronal
35100838|T121|Endronax
35100837|T121|Endrostan
35100836|T121|Endrox
35100835|T121|Epidexone
35100834|T121|Epidrone
35100833|T121|Epizolone
35100832|T121|Erbanfol
35100831|T121|Erladexone
35100830|T121|Ermethasone
35100829|T121|Eroprim
35100828|T121|Erotrim
35100827|T121|Erphatrim
35100826|T121|Esbesul
35100825|T121|Escoprim
35100824|T121|Espasevit
35100823|T121|Espectrin
35100822|T121|Espectroprima
35100821|T121|Estroquin
35100820|T121|ETA Cortilen
35100819|T121|Etason
35100818|T121|Ethitrim
35100817|T121|Eucalen
35100816|T121|Euromethasone
35100815|T121|Eurotrim
35100814|T121|Eusaprim
35100813|T121|Eutrim
35100812|T121|Exazol
35100811|T121|Excelin
35100810|T121|Exemestane and Tucidinostat
35100809|T121|Fabubac
35100808|T121|Fada Dexametasona
35100807|T121|Fadametasona
35100806|T121|Fakzol
35100805|T121|Falprim
35100804|T121|Fameprim
35100803|T121|Faridexon
35100802|T121|Farin
35100801|T121|Fastovorin
35100800|T121|Fauldleuco
35100799|T121|Fayining
35100798|T121|Fectrim
35100797|T121|Fedimed
35100796|T121|Fedolen
35100795|T121|Fentul
35100794|T121|Ferbon
35100793|T121|Ferevan
35100792|T121|Fericard
35100791|T121|Feron
35100790|T121|Fexadron
35100789|T121|Fiblaferon
35100788|T121|Finaber
35100787|T121|Findeclin
35100786|T121|Finnferon-Alpha
35100785|T121|Finoxi
35100784|T121|Firmofos
35100783|T121|Fisat
35101450|T121|Fixopan
35101449|T121|Flatran
35101448|T121|Flocot
35101447|T121|Fluril
35101446|T121|Folaren
35101445|T121|Folaxin
35101444|T121|Folend
35101443|T121|Foli Cell
35101442|T121|Foliben
35101441|T121|Folidan
35101440|T121|Folidar
35101439|T121|Foliment
35101438|T121|Folinac
35101437|T121|Folinato
35101436|T121|Folinfabra
35101435|T121|Folinoral
35101434|T121|Folinoxan
35101433|T121|Folinvit
35101432|T121|Foliplus
35101431|T121|Folmigor
35101430|T121|Forcrim
35101429|T121|Forenmax
35101428|T121|Fortecortin
35101427|T121|Forteprim
35101426|T121|Fosaalen
35101425|T121|Fosalan
35101424|T121|Fosalen
35101423|T121|Fosalong
35101422|T121|Fosamac
35101421|T121|Fosamax
35101420|T121|Fosanet
35101419|T121|Fosaqueen
35101418|T121|Fosavance
35101417|T121|Fosfalen
35101416|T121|Fosfato Dissodico Dexametasona
35101415|T121|Fosfidex
35101414|T121|Fosfoplus
35101413|T121|Fosmin
35101412|T121|Fostepor
35101411|T121|Fosval
35101410|T121|Frazon
35101409|T121|Frone
35101408|T121|Gamactrin
35101407|T121|Gammacorten
35101406|T121|Gatrima
35101405|T121|Gemisona
35101404|T121|Genalen
35101403|T121|Genalmen
35101402|T121|Genoctrin
35101401|T121|Genoxzole
35101400|T121|Gentrim
35101399|T121|Genzaprim
35101398|T121|Gerical
35101397|T121|Getrim
35101396|T121|Glendan
35101395|T121|Globaxol
35101394|T121|Glymesason
35101393|T121|Gobens Trim
35101392|T121|Graprima
35101391|T121|Grathazon
35101390|T121|Groseptol
35101389|T121|Gunametrim
35101388|T121|Gynodron
35101387|T121|Haemofarin
35101386|T121|Haloxan
35101385|T121|Hatrix
35101384|T121|Heberon Alfa R
35101383|T121|Helmine
35101382|T121|Helveprim
35101381|T121|Herixina
35101380|T121|Hexadecadrol
35101379|T121|Hexadrol
35101378|T121|Hexaprim
35101377|T121|Hexilon
35101376|T121|HI-Methasone
35101375|T121|Hicot
35101374|T121|Holadren
35101373|T121|Holoxan
35101372|T121|Holoxane
35101371|T121|Hopamethasone
42542448|T121|HPV-positive Oropharyngeal cancer
35101370|T121|Hufacid
35101369|T121|Huma-Trimel
35101368|T121|Humoferon
35101367|T121|Ibrunib
35101366|T121|Ibrutix
35101365|T121|Ibtrim
35101364|T121|Idizone
35101363|T121|Ifavor
35101362|T121|Ifex
35101361|T121|IFN Alpha
35101360|T121|IFO Cell
35101359|T121|Ifocris
35101358|T121|Ifolem
35101357|T121|Ifomida
35101356|T121|Ifomide
35101355|T121|Ifos
35101354|T121|Ifosfamida
35101353|T121|Ifoxan
35101352|T121|IFX
35101351|T121|Imatinib, Vincristine, Prednisone
35101350|T121|Imcotran
35101349|T121|Imexim
35101348|T121|Imufor
35101347|T121|Imukin
35101346|T121|Inatrim
35101345|T121|Indexon
35101344|T121|Indrol
35101343|T121|INF
35101342|T121|Infatrim
35101341|T121|Infectran
35101340|T121|Infectrim
35101339|T121|Infectrin
35101338|T121|Inferax
35101337|T121|Infergen
35101336|T121|Infesin
35101335|T121|Injectrax
35101334|T121|Inmutag
35101333|T121|Insetron
35101332|T121|Interfero
35101331|T121|Interferon Alfanative
35101330|T121|Interferon Human
35101329|T121|Interferon Leucocyticum
35101328|T121|Interferon Lymphoblastoid
35101327|T121|Interferonum Leucocyticum
35101326|T121|Interval debulking surgery
35101325|T121|Inthesa-5
35101324|T121|Intidrol
35101323|T121|Intrafort
35101322|T121|Introcin
35101321|T121|Invomit
35101320|T121|Ipamide
35101319|T121|Irgagen
35101318|T121|Irinomedac
35101317|T121|Irzamethazone
35101316|T121|Isodexam
35101315|T121|Isophosphamide
35101314|T121|Isoprim
35101313|T121|Isopto
35101312|T121|Isotretinoin and Dinutuximab
35101311|T121|Isotrim
35101310|T121|Isovorin
35101309|T121|Isoxan
35101308|T121|Ivepred
35101307|T121|Izofran
35101306|T121|Jantoven
35101305|T121|Japtrim
35101304|T121|Jasotrim
35101303|T121|Jenamoxazol
35101302|T121|Jestrim
35101301|T121|Justeprim
35101300|T121|K.B.famate
35101299|T121|Kaarmepakkaus
35101298|T121|Kaftrim
35101297|T121|Kalciumfolinat Perivita
35101296|T121|Kalmethasone
35101295|T121|Kalsiumfolinat
35101294|T121|Kanadex
35101293|T121|Kathrex
35101292|T121|Katrim
35101291|T121|Kaytran
35101290|T121|Keflex
35101289|T121|Kemocid
35101288|T121|Kemoprim
35101287|T121|Kentricid
35100782|T121|Kepinol
35100781|T121|Kepivance
35100780|T121|Kindoprim
35100779|T121|KO-Kure
35100778|T121|Kodolo
35100777|T121|Kombina
35100776|T121|Kosa
35100775|T121|Kotazol
35100774|T121|Kotrimoksazol
35100773|T121|Kovar
35100772|T121|Kovintong
35100771|T121|Krobactrol
35100770|T121|Kunyrin
35100769|T121|L-Trim
35100768|T121|Lacreozole
35100767|T121|Lafedam
35100766|T121|Lagatrim
35100765|T121|Lameson
35100764|T121|Lanadexon
35100763|T121|Landrolen
35100762|T121|Lapikot
35100761|T121|Laratrim
35100760|T121|Laroferon
35100759|T121|Larprim
35100758|T121|Lastrim
35100757|T121|Latran
35100756|T121|Lawarin
35100755|T121|Lederfolat
35100754|T121|Lederfolin
35100753|T121|Lederfoline
35100688|T121|Ledervorin
35100687|T121|Legifol
35100686|T121|Lemod
35100685|T121|Lendronal
35100684|T121|Leodrin
35100683|T121|Leotrim
35100682|T121|Leprim
35100681|T121|Lescot
35100680|T121|Lesol
35100679|T121|Letus
35100678|T121|Leucocalcin
35100677|T121|Leuconolver
35100676|T121|Leucovorin
35100675|T121|Leucovorina
35100674|T121|Leucovorine
35100673|T121|Leukeran
35100672|T121|Leukovorin
35100671|T121|Lexcomet
35100670|T121|Lexxema
35100669|T121|Licoson
35100668|T121|Lictora
35100667|T121|Lifactrin
35100666|T121|Lifzol
35100665|T121|Limethason
35100664|T121|Lindron
35100663|T121|Linfoxan
35100662|T121|Lipotalon
35100661|T121|Lisaprin
35100660|T121|Lisoderme
35100659|T121|Litrim
35100658|T121|Lobact
35100657|T121|Lodex
35100656|T121|Lodexa
35100655|T121|Lokalison-F
35100654|T121|Lokar
35100653|T121|Lomustine, Temozolomide, RT
35100653|T121|Lomustine, Temozolomide, Radiation Therapy
35100652|T121|Longasal
35100651|T121|Lormine
35100650|T121|Loverine
35100649|T121|Lovorin
35100648|T121|Lucibru
35100647|T121|Lupectrin
35100646|T121|Lupidexa
35100645|T121|Lusaprim
35100644|T121|Luxazone
35100643|T121|Lykaprim
35100642|T121|M-Moxa
35100641|T121|M-Prednihexal
35100640|T121|M-Trim
35100639|T121|Macdafen
35100638|T121|Macprim
35100637|T121|Macromed
35100636|T121|Mactran
35100635|T121|Madroxin
35100634|T121|Maforan
35100633|T121|Maktrim
35100632|T121|Maradex
35100631|T121|Marfarin
35100630|T121|Marivanil
35100629|T121|Marivarin
35100628|T121|Martiprim
35100627|T121|Marvil
35100626|T121|Maxaprim
35100625|T121|Maxibone
35100624|T121|Maxidex
35100623|T121|Maxiprim
35100622|T121|Maxitrin
35100621|T121|Maxol
35100620|T121|Maxtrim
35100619|T121|Maxzol
35100618|T121|Mazatrim
35100617|T121|MBVP
35100617|T121|Methotrexate, BCNU (Carmustine), Vumon (Teniposide), Prednisone
35100616|T121|Mebryn
35100615|T121|Mecoxon
35100614|T121|Medason
35100613|T121|Medcotrim
35100612|T121|Medesone
35100611|T121|Medexasone
35100610|T121|Mediamethasone
35100609|T121|Medicofolin
35100608|T121|Medidex
35100607|T121|Medifolin
35100606|T121|Mediprim
35100605|T121|Medirona
35100604|T121|Medisolu
35100603|T121|Meditran
35100602|T121|Meditrim
35100601|T121|Medixon
35100600|T121|Medlin
35100599|T121|Medlone
35100598|T121|Mednin
35100597|T121|Medralone
35100596|T121|Medrate
35100595|T121|Medrol
35100594|T121|Medrone
35100593|T121|Medsavorina
35100592|T121|Medtrim
35100591|T121|Megabroncoflam
35100590|T121|Megacort
35100589|T121|Megadex
35100588|T121|Megaset
35100587|T121|Megatrim
35100586|T121|Melon
35100585|T121|Melone
35100584|T121|Menisolon
35100583|T121|Menisone
35100582|T121|Mephameson
35100581|T121|Mephamesona
35100580|T121|Mephamesone
35100579|T121|Mephamesone-4
35100578|T121|Mepredron
35100577|T121|Meprim
35100576|T121|Meprolone Unipak
35100575|T121|Meproson
35100574|T121|Meprotrin
35100573|T121|Mepsolone
35100572|T121|Mepson
35100571|T121|Meradexon
35100570|T121|Merideca
35100569|T121|Mesadoron
35100568|T121|Mesolone
35100567|T121|Mesurin
35100566|T121|Metalexina
35100565|T121|Metasolon
35100564|T121|Metax
35100563|T121|Metaxon
35100562|T121|Metcort
35100561|T121|Methaderm
35100560|T121|Methapred
35100559|T121|Methasone
35100558|T121|Methisol
35100557|T121|Methoprim
35100556|T121|Methotrin
35100555|T121|Methybon
35100554|T121|Methylon
35100553|T121|Methylone
35100552|T121|Methylprednis
35100551|T121|Methylprednisolon
35100550|T121|Methylprednisolonum
35100549|T121|Methyran
35100548|T121|Meticort
35100547|T121|Metidrol
35100546|T121|Metilbetasone
35100545|T121|Metilprednisolona
35100544|T121|Metilprednizolon-H
35100543|T121|Metipred
35100542|T121|Metisone
35100541|T121|Metoprim
35100540|T121|Metoprin
35100539|T121|Metoxiprim
35100538|T121|Metrim
35100537|T121|Metxaprim
35100536|T121|Metycortin
35100535|T121|Metypred
35100534|T121|Metypresol
35100533|T121|Metysolon
35100532|T121|Mexaprim
35100531|T121|Mexasone
35100530|T121|Mexaton
35100529|T121|Mexazole
35100528|T121|Mezenol
35100527|T121|Micinovo
35100526|T121|Micogyl
35100525|T121|Microbid
35100524|T121|Microcetim
35100523|T121|Microdyn
35100522|T121|Microsupos Amigdalar
35100521|T121|Microtrim
35100520|T121|Migradexan
35100519|T121|Mikotrim
35100518|T121|Mikrosid
35100517|T121|Millicorten
35100516|T121|Minidex
35100515|T121|Minusorb
35100514|T121|Miratrim
35100513|T121|Mitasone
35100512|T121|Mitoxana
35100511|T121|Modifical
35100510|T121|Molacort
35100509|T121|Moly
35100508|T121|Monkast
35100507|T121|Montair
35100506|T121|Mortin
35100505|T121|Moxadden
35100504|T121|Moxalas
35100503|T121|Moxatrim
35101070|T121|Moxzole
35101069|T121|Mukadryl
35101068|T121|Multiferon
35101067|T121|Mycidex
35101066|T121|Mycostatin
35101065|T121|Myctrim
35101064|T121|Naftran
35101063|T121|Namalvin
35101062|T121|Napatrim
35101061|T121|Narfoz
35101060|T121|Nausedron
35101059|T121|Nautah
35101058|T121|Navatrim
35101057|T121|Necorzole
35101056|T121|NEO-Drol
35101055|T121|Neodex
35101054|T121|Neofolin
35101053|T121|Neomit
35101052|T121|Neoset
35101051|T121|Neotrim
35101050|T121|Netocur
35101049|T121|Neuroprim
35101048|T121|Nexadron
35101047|T121|Nichospor
35101046|T121|Nicotrim
35101045|T121|Nilium
35101044|T121|Nirypan
35101043|T121|Nodevex
35101042|T121|Nodilon
35101041|T121|Nopil
35101040|T121|Norisep
35101039|T121|Nortrim
35101038|T121|Nortrime
35101037|T121|Notrim
35101036|T121|Notrime
35101035|T121|Novactil
35101034|T121|Novidrine
35101033|T121|Novotrim Plus
35101032|T121|Novotrimel
35101031|T121|Novotrimox
35101030|T121|Novozole
35101029|T121|Nucotrim
35101028|T121|Nufadex M
35101027|T121|Nufaprim
35101026|T121|Nuruzole
35101025|T121|Nuset
35101024|T121|Nyrin
35101023|T121|Nystatin
35101022|T121|O Folin
35101021|T121|O.N.D.
35101020|T121|Ocedran
35101019|T121|Octil-S
35101018|T121|Octran
35101017|T121|Octrim
35101016|T121|Ocudex
35101015|T121|Odanex
35101014|T121|Odanse
35101013|T121|Oecotrim
35101012|T121|Oftadek
35101011|T121|Oftadex
35101010|T121|OIF
35101009|T121|Okatrim
35101008|T121|Omedexon
35101007|T121|Omegtrim
35101006|T121|Ometic
35101005|T121|Omnatrim
35101004|T121|Omsat
35101003|T121|Omstron
35101002|T121|Onadron
35101001|T121|Onaset
35101000|T121|Onclast
35100999|T121|Oncotor
35100998|T121|Oncovin
35100997|T121|Onda
35100996|T121|Ondace
35100995|T121|Ondan
35100994|T121|Ondanles
35100993|T121|Ondansetron-Z
35100992|T121|Ondant
35100991|T121|Ondaren
35100990|T121|Ondasetron
35100989|T121|Ondatie
35100988|T121|Ondavell
35100987|T121|Ondem
35100986|T121|Ondemet
35100985|T121|Onetrim
35100984|T121|Onfran
35100983|T121|Onilat
35100982|T121|Onsat
35100981|T121|Onseran
35100980|T121|Onset
35100979|T121|Onsetron
35100978|T121|Onsett
35100977|T121|Onsia
35100976|T121|Ontrax
35100975|T121|Onzod
35100974|T121|Ophth-DEX
35100973|T121|Ophthasona
35100972|T121|Opticort
35100971|T121|Optune
35100970|T121|Oradin
35100969|T121|Orazone
35100502|T121|Orbak
35100501|T121|Ordex
35100500|T121|Orfarin
35100499|T121|Orgadrone
35100498|T121|Orgastran
35100497|T121|Oribact
35100496|T121|Ormoprim
35100495|T121|Orthonate
35100494|T121|Osalen
35100493|T121|Osaston
35100492|T121|Osdronat
35100491|T121|Oseolen
35100490|T121|Oseomax
35100489|T121|Oseotal
35100488|T121|Oseotenk
35100487|T121|Osetron
35100486|T121|Osficar
35100485|T121|Osfolate
35100484|T121|Osfolato
35100483|T121|Oslene
35100482|T121|Ossifix
35100481|T121|Ossomax
35100480|T121|Ostasyn
35100479|T121|Ostat
35100478|T121|Ostel
35100477|T121|Ostemax Comfort
35100476|T121|Ostenan
35100475|T121|Osteobon
35100474|T121|Osteodur
35100473|T121|Osteofar
35100472|T121|Osteofel
35100471|T121|Osteofene
35100470|T121|Osteofos
35100469|T121|Osteofose
35100468|T121|Osteomax
35100467|T121|Osteomed
35100466|T121|Osteomel
35100465|T121|Osteomepha
35100464|T121|Osteomix
35100463|T121|Osteonato
35100462|T121|Osteoral
35100461|T121|Osteotec
35100460|T121|Osteotrat
35100459|T121|Ostex
35100458|T121|Ostolek
35100457|T121|Ostonat
35100456|T121|Ostrin Forte
35100455|T121|Otobrol
35100454|T121|Otrim
35100453|T121|Ottoprim
35100452|T121|Oxaprim
35100451|T121|Oxtalen
35100450|T121|Pakzole
35100449|T121|rhKGF
35100449|T121|Palifermin
35100448|T121|Pantrim
35100447|T121|Panwarfin
35100446|T121|Panwarfine
35100445|T121|Patrim
35100444|T121|Pegfilgrastim-cbqv
35100443|T121|Pehatrim
35100442|T121|Penatone
35100441|T121|Penetrin
35100440|T121|Penicillin
35100439|T121|Penicillin V
35100438|T121|Penodex
35100437|T121|Pentrin
35100436|T121|Penzole
35100435|T121|Perfolate
35100434|T121|Periset
35100433|T121|Peyrone's Chloride
35100432|T121|Peyrone's Salt
35100431|T121|Phadilon
35100430|T121|Pharmatrim
35100429|T121|Pharmazol
35100428|T121|Phartex
35100427|T121|Phenodex
35100426|T121|Phostarac
35100425|T121|Pidexon
42542449|T121|PIK3CA-mutated Breast cancer
35100424|T121|Piqray
35100423|T121|Pisatrina
35100422|T121|Plastistil
35100421|T121|Platinex
35100420|T121|Plavex
35100419|T121|Plenair
35100418|T121|Plidexa
35100417|T121|Plurisul
35100416|T121|DCDS4501A
35100416|T121|polatuzumab vedotin-piiq
35100416|T121|Polatuzumab vedotin
35100415|T121|Polibatrin
35100414|T121|Politrim
35100413|T121|Polivy
35100412|T121|Polyferon
35100411|T121|Polytran
35100410|T121|Poris
35100409|T121|Porosal
35100408|T121|Porosin
35100407|T121|Predisol
35100406|T121|Predmetil
35100405|T121|Predni M
35100404|T121|Predni-M-Tablinen
35100403|T121|Prednilem
35100402|T121|Prednol
35100401|T121|Prednol L
35100400|T121|Prednovare
35100399|T121|Prednox
35100398|T121|Prefolic
35100397|T121|Pretilon
35100396|T121|Prevax
35100395|T121|Pribac
35100394|T121|Pridol
35100393|T121|Primadex
35100392|T121|Primasul
35100391|T121|Primasulf
35100390|T121|Primatrim
35100389|T121|Primavon
35100388|T121|Primazol
35100387|T121|Primazole
35100386|T121|Primotren
35100385|T121|Primox
35100384|T121|Primsulfon
35100383|T121|Primzole
35100382|T121|Prodexon
35100381|T121|Promedrol
35100380|T121|Protrin
35100379|T121|Pulkrin
35100378|T121|Purbac
35100377|T121|Pyderma
35100376|T121|Pyradexon
35100375|T121|Qiftrim
35100374|T121|Qiftrin
35100373|T121|Quimio-PED
35100372|T121|Quimiofran
35100371|T121|Quisulyn
35100370|T121|Radilem
35100369|T121|Ralenost
35100368|T121|Rally-A
35100367|T121|Rancotrim
35100366|T121|Randexa
35100365|T121|Rasat
35100364|T121|Raseptol
35100363|T121|Ratrim
35100362|T121|ravulizumab-cwvz
35100362|T121|ALXN1210
35100362|T121|Ravulizumab
35100361|T121|Ravulizumab monotherapy
35100360|T121|Realdiron
35100359|T121|Recalfe
35100358|T121|Recovorin
35100357|T121|Redexon
35100356|T121|Rednisone
35100355|T121|Regenesis
35100354|T121|Regtin
35100353|T121|Rekostin
35100352|T121|Rematrim
35100351|T121|Renatrim
35100350|T121|Reotan
35100349|T121|Rescuvolin
35100348|T121|Resfolin
35100347|T121|Resprim
35100346|T121|Restofos
35100345|T121|Retrim
35100344|T121|Reusan
35100343|T121|Reventa
35100342|T121|Rexaprim
35100341|T121|Ribatrim
35100340|T121|Ribofolin
35100339|T121|Rimazole
35100338|T121|Rimezone
35100337|T121|Rivoprim
35100336|T121|Rizol
35100335|T121|Roceron-A
35100334|T121|Rocolone
35100333|T121|Rolprim
35100332|T121|Romax
35100331|T121|Romesa
35100330|T121|Ronic
35100329|T121|Rontafor
35100328|T121|Roubac
35100327|T121|Roximeth
35100326|T121|Roxtrim
35100325|T121|Roytrin
35100324|T121|Rumaxoi
35100323|T121|Rupedex
35100322|T121|Salgatran
35100321|T121|Salon H9C
35100320|T121|Saltrim
35100319|T121|Samofaron
35100318|T121|Sanexon
35100317|T121|Sanifolin
35100316|T121|Sanprima
35100315|T121|Santeson
35100314|T121|Saptrim
35100313|T121|Satrim
35100312|T121|Sawasone
35100311|T121|Sbpa Trimeth Smeth
35100310|T121|Scandexon
35100309|T121|Scribcin
35100308|T121|Seematrim
35100307|T121|Seftrim
35100306|T121|Selectrin
35100305|T121|Selftison
35100304|T121|Selinexor and Dexamethasone (Sd)
35100304|T121|Sd
35100304|T121|Selinexor and low-dose dexamethasone
35100303|T121|Semozol
35100302|T121|Sepiran
35100301|T121|Sepmax
35100300|T121|Septabid
35100299|T121|Septazol
35100298|T121|Septazole
35100297|T121|Septerin
35100296|T121|Septinix
35100295|T121|Septiolan
35100294|T121|Septocid R +
35100293|T121|Septoprin
35100292|T121|Septra
35100291|T121|Septran
35100290|T121|Septrin Paediatric
35100289|T121|Septrin-S
35100288|T121|Servitrim
35100287|T121|Seton
35100752|T121|Setronax
35100751|T121|Setronon
35100750|T121|Shirodex
35100749|T121|Shuayan
35100748|T121|Sigaprim
35100747|T121|Sigatrim
35100746|T121|Silidral
35100745|T121|Silpin
35100744|T121|Siltran
35100743|T121|Simarc
35100742|T121|Sinatrim
35100741|T121|Sinersul
35100740|T121|Sinfract
35100739|T121|Singulair
35100738|T121|Sinotrim
35100737|T121|Sisoprim
35100736|T121|Sistrim
35100735|T121|Sitrim
35100734|T121|Skytrin
35100733|T121|Smartrim
35100732|T121|Smile
35100731|T121|SOL-Melcort
35100730|T121|Solcort
35100729|T121|Soldesam
35100728|T121|Soldesanil
35100727|T121|Soldex
35100726|T121|Solocort-ACT
35100725|T121|Solomet
35100724|T121|Soltrim
35100723|T121|Solu Moderin
35100722|T121|Soludecadron
35100721|T121|Solumedrol
35100720|T121|Solupen
35100719|T121|Somelon
35100718|T121|Somerol
35100717|T121|Sonexa
35100716|T121|Sopran
35100715|T121|Soptrim
35100714|T121|Sosetran
35100713|T121|SP Cordexa
35100712|T121|Spectrem
35100711|T121|Spectrim
35100710|T121|Spersadex
35100709|T121|Spondy-Dexa
35100708|T121|Stan
35100707|T121|Stedex
35100706|T121|Stenirol
35100705|T121|Steralol
35100704|T121|Sterasone
35100703|T121|Steron
35100702|T121|Stopan
35100701|T121|Strim
35100700|T121|Strontium-89
35100699|T121|Succimed
35100698|T121|Suftrex
35100697|T121|Sulbacta
35100696|T121|Sulfagrand
35100695|T121|Sulfamer
35100694|T121|Sulfamet
35100693|T121|Sulfamethoprim
35100692|T121|Sulfametoxazol
35100691|T121|Sulfaprim
35100690|T121|Sulfarim
35100689|T121|Sulfatalpin
35100286|T121|Sulfaton
35100285|T121|Sulfatrim
35100284|T121|Sulfatropim
35100283|T121|Sulfawal-T
35100282|T121|Sulfinam
35100281|T121|Sulfoid Trimetho
35100280|T121|Sulfometh
35100279|T121|Sulfonamide
35100278|T121|Sulfort
35100277|T121|Sulfotrim
35100276|T121|Sulfotrimin
35100275|T121|Sulftran
35100274|T121|Sulgotri
35100273|T121|Sulotrim
35100272|T121|Sulphaprim
35100271|T121|Sulphathoprim
35100270|T121|Sulphatran
35100269|T121|Sulphatrim
35100268|T121|Sulphax
35100267|T121|Sulphytrim Forte
35100266|T121|Sulprim
35100265|T121|Sulprimed
35100264|T121|Sultase
35100263|T121|Sulthrim
35100262|T121|Sultiprim
35100261|T121|Sultorim
35100260|T121|Sultra
35100259|T121|Sultrex
35100258|T121|Sultrim
35100257|T121|Sultrima
35100256|T121|Sultrimmix
35100255|T121|Sultrivon-F
35100254|T121|Sultropim
35100253|T121|Sumetoprim
35100252|T121|Sumetrolim
35100251|T121|Sumetrolin
35100250|T121|Sumiferon
35100249|T121|Sumitran
35100248|T121|Suntrim
35100247|T121|Superprednol
35100246|T121|Supertendin-Depot N
35100245|T121|Supim
35100244|T121|Supracombin
35100243|T121|Suprason
35100242|T121|Suprasulf
35100241|T121|Suprax
35100240|T121|Supresol
35100239|T121|Suprex
35100238|T121|Supribac
35100237|T121|Suprim
35100236|T121|Suprimass
35100235|T121|Suprin
35100234|T121|Suptrex
35100233|T121|Suptrim
35100232|T121|Surodex
35100231|T121|Sutaprim
35100230|T121|Sutrim
35100229|T121|Sutrisan
35100228|T121|Suxprim
35100227|T121|Sydencort
35100226|T121|Syltrifil
35100225|T121|Synac
35100224|T121|Synastat
35100223|T121|Synbac
35100222|T121|Synco-Smzt
35100221|T121|Syndal
35100220|T121|Syndexa
35100219|T121|Synermed
35100218|T121|Synerzole
35100217|T121|Synetra
35100216|T121|Synostep
35100215|T121|Synotrim
35100214|T121|Syntoprim
35100213|T121|System
35100212|T121|Tabrol
35100211|T121|Tagremin
35100210|T121|Tavesona
35100209|T121|Teanlang
35100208|T121|Tecnovorin
35100207|T121|Tedicumar
35100206|T121|Teikason Nidek
35100205|T121|Teiroc
35100204|T121|Tekuron
35100203|T121|Teof
35100202|T121|Terasulf
35100201|T121|Terbosulfa
35100200|T121|Terost
35100199|T121|Teutrin
35100198|T121|Tevalen
35100197|T121|Tevanate
35100196|T121|Theraprim
35100195|T121|Therasept
35100194|T121|Theratrim
35100193|T121|Thilodex
35100192|T121|Thilodexine
35100191|T121|Thimelon
35100190|T121|Thoprim
35100189|T121|Thriazol
35100188|T121|Thymitaq
35100187|T121|Tibolene
35100186|T121|Tibone
35100185|T121|Tilios
35100184|T121|Tonofolin
35100183|T121|Torisel
35100182|T121|Torrid
35100181|T121|Totocortin
35100180|T121|Tprim
35100178|T121|Trelibec
35100177|T121|Trib
35100176|T121|Tricban
35100175|T121|Tricomox
35100174|T121|Tricot
35100173|T121|Trifides
35100172|T121|Triforam
35100171|T121|Trihexal
35100170|T121|Trim
35100169|T121|Trima
35100168|T121|Trimaxazole
35100167|T121|Trimel
35100166|T121|Trimephar
35100165|T121|Trimeran
35100164|T121|Trimerazin
35100163|T121|Trimeril
35100162|T121|Trimesol
35100161|T121|Trimesul
35100160|T121|Trimesulf
35100159|T121|Trimeta
35100158|T121|Trimethox
35100157|T121|Trimetoger
35100156|T121|Trimetop Duplo
35100155|T121|Trimetotal
35100154|T121|Trimetox
35100153|T121|Trimetrin
35100152|T121|Trimetsol
35100151|T121|Trimexasol
35100150|T121|Trimexazol
35100149|T121|Trimexazole
35100148|T121|Trimexole-F
35100147|T121|Trimezol
35100146|T121|Trimezole
35100145|T121|Trimfasul
35100144|T121|Trimidar M
35100143|T121|Triminex
35100142|T121|Trimocom
35100141|T121|Trimoks
35100140|T121|Trimosul
35100139|T121|Trimosulfa
35100138|T121|Trimoxavin
35100137|T121|Trimoxazol
35100179|T121|Trimoxazole-BC
35100136|T121|Trimoxin
35100135|T121|Trimoxis
35100134|T121|Trimoxsul
35100133|T121|Trimozol
35100132|T121|Trimsul
35100131|T121|Trimzol
35100130|T121|Triphimox
35100129|T121|Tripur
35100128|T121|Trisep
35100127|T121|Trisfides
35100126|T121|Trisolak Forte
35100125|T121|Trisolvat
35100124|T121|Trisul
35100123|T121|Trisulcom
35100122|T121|Trisulfa
35100121|T121|Trisulfose
35100120|T121|Trisuprim
35100119|T121|Trisural
35100118|T121|Tritenk
35100117|T121|Tritosul
35100116|T121|Trixazol
35100115|T121|Trixzol
35100114|T121|Trizole
35100113|T121|Tronoxal
35100112|T121|Tropidrol
35100111|T121|Trorix
35100110|T121|Tryseptolum
35100109|T121|Tuttozem N
35100108|T121|Tytrim
35100107|T121|U-Prin
35100106|T121|Ucalon
35100105|T121|Udicort
35100104|T121|Ulfaprim
35100103|T121|Ultomiris
35100102|T121|Ultrasept
35100101|T121|Ultrazole
35100100|T121|Ultrim
35100099|T121|Unidex
35100098|T121|Unidexa
35100097|T121|Unimedrol
35100096|T121|Unisone
35100095|T121|Unitran
35100094|T121|Uprina
35100093|T121|Urbason
35100092|T121|Urethrax
35100091|T121|Urodown
35100090|T121|Uroplus DS
35100089|T121|Urtium
35100088|T121|Utrin
35100087|T121|Vanderm
35100086|T121|Varfarins
35100085|T121|Varfine
35100084|T121|Venetoclax and Obinutuzumab
35100084|T121|VG
35100084|T121|VO
35100084|T121|GVE
35100084|T121|Venetoclax and Gazyva (Obinutuzumab)
35100084|T121|Gazyva (Obinutuzumab) and VEnetoclax
35100083|T121|Veravorin
35100082|T121|Versatrim
35100081|T121|Ves-ATRA
35100080|T121|Vesanoid
35100079|T121|Virin
35100078|T121|Visualin
35100077|T121|Visumetazone
35100076|T121|Voalla
35100075|T121|Vomceran
35100074|T121|Vomiban
35100073|T121|Vomigo
35100072|T121|Vomikind
35100071|T121|Vomiset
35100070|T121|Vomitron
35100069|T121|Vomiz
35100068|T121|Vonau
35100067|T121|Vorina
35100066|T121|Voroste
35100065|T121|Waran
35100064|T121|Warf
35100063|T121|Warfa
35100062|T121|Warfant
35100061|T121|Warfar
35100060|T121|Warfarex
35100059|T121|Warfil
35100058|T121|Warfilone
35100057|T121|Warfin
35100056|T121|Warin
35100055|T121|Warlin
35100054|T121|Warnerin
35100053|T121|Weiditrin
35100052|T121|Wellcovorin
35100051|T121|Wellferon
35100050|T121|Werifrin
35100049|T121|Wiatrim
35100048|T121|Wiltran
35100047|T121|Windex
35100046|T121|Wymesone
35100045|T121|Wypal
35100044|T121|X-Trim
35100043|T121|XA-Zole
35100042|T121|Xasone
35100041|T121|Xazotrim
35100040|T121|Xepaprim
35100039|T121|Xerazole
35100038|T121|Xeroprim
35100037|T121|Xine
35100036|T121|Xpovio
35100035|T121|Yatrox
35100034|T121|Yekaprim
35100033|T121|Yumerole
35100032|T121|Zactron
35100031|T121|Zalucs
35100030|T121|Zamboprim
35100029|T121|Zantran
35100028|T121|Zantron
35100027|T121|Zapron
35100026|T121|Zaxol
35100025|T121|Zecatrim
35100024|T121|Zecaxon
35100023|T121|Zemitron
35100022|T121|Zenos
35100021|T121|Zeptra
35100020|T121|Zerrprim
35100019|T121|Zirabev
35100018|T121|Zofer
35100017|T121|Zofran
35100016|T121|Zofran ODT
35100015|T121|Zofron
35100014|T121|Zolebid
35100013|T121|Zolmed
35100012|T121|Zoltem
35100011|T121|Zoltrijem
35100010|T121|Zoltrim
35100009|T121|Zonax
35100008|T121|Zondan
35100007|T121|Zophost
35100006|T121|Zophren
35100005|T121|Zudan
35100004|T121|Zultrop
35100003|T121|Zydexa
35100002|T121|Zyofolin
35100001|T121|Zytofolin
912262|T121|Boniva
