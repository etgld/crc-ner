000|T121|TC
000|T121|Taxotere
000|T121|Cytoxan