000|T121|chemotherapy
000|T121|chemotherapies
000|T121|chemo
000|T121|chemotherapeutic
000|T121|cytoxan
000|T121|taxotere
000|T121|tamoxifen
000|T121|tc